
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"41",x"7f",x"7f",x"00"),
     1 => (x"01",x"00",x"00",x"41"),
     2 => (x"18",x"0c",x"06",x"03"),
     3 => (x"00",x"40",x"60",x"30"),
     4 => (x"7f",x"41",x"41",x"00"),
     5 => (x"08",x"00",x"00",x"7f"),
     6 => (x"06",x"03",x"06",x"0c"),
     7 => (x"80",x"00",x"08",x"0c"),
     8 => (x"80",x"80",x"80",x"80"),
     9 => (x"00",x"00",x"80",x"80"),
    10 => (x"07",x"03",x"00",x"00"),
    11 => (x"00",x"00",x"00",x"04"),
    12 => (x"54",x"54",x"74",x"20"),
    13 => (x"00",x"00",x"78",x"7c"),
    14 => (x"44",x"44",x"7f",x"7f"),
    15 => (x"00",x"00",x"38",x"7c"),
    16 => (x"44",x"44",x"7c",x"38"),
    17 => (x"00",x"00",x"00",x"44"),
    18 => (x"44",x"44",x"7c",x"38"),
    19 => (x"00",x"00",x"7f",x"7f"),
    20 => (x"54",x"54",x"7c",x"38"),
    21 => (x"00",x"00",x"18",x"5c"),
    22 => (x"05",x"7f",x"7e",x"04"),
    23 => (x"00",x"00",x"00",x"05"),
    24 => (x"a4",x"a4",x"bc",x"18"),
    25 => (x"00",x"00",x"7c",x"fc"),
    26 => (x"04",x"04",x"7f",x"7f"),
    27 => (x"00",x"00",x"78",x"7c"),
    28 => (x"7d",x"3d",x"00",x"00"),
    29 => (x"00",x"00",x"00",x"40"),
    30 => (x"fd",x"80",x"80",x"80"),
    31 => (x"00",x"00",x"00",x"7d"),
    32 => (x"38",x"10",x"7f",x"7f"),
    33 => (x"00",x"00",x"44",x"6c"),
    34 => (x"7f",x"3f",x"00",x"00"),
    35 => (x"7c",x"00",x"00",x"40"),
    36 => (x"0c",x"18",x"0c",x"7c"),
    37 => (x"00",x"00",x"78",x"7c"),
    38 => (x"04",x"04",x"7c",x"7c"),
    39 => (x"00",x"00",x"78",x"7c"),
    40 => (x"44",x"44",x"7c",x"38"),
    41 => (x"00",x"00",x"38",x"7c"),
    42 => (x"24",x"24",x"fc",x"fc"),
    43 => (x"00",x"00",x"18",x"3c"),
    44 => (x"24",x"24",x"3c",x"18"),
    45 => (x"00",x"00",x"fc",x"fc"),
    46 => (x"04",x"04",x"7c",x"7c"),
    47 => (x"00",x"00",x"08",x"0c"),
    48 => (x"54",x"54",x"5c",x"48"),
    49 => (x"00",x"00",x"20",x"74"),
    50 => (x"44",x"7f",x"3f",x"04"),
    51 => (x"00",x"00",x"00",x"44"),
    52 => (x"40",x"40",x"7c",x"3c"),
    53 => (x"00",x"00",x"7c",x"7c"),
    54 => (x"60",x"60",x"3c",x"1c"),
    55 => (x"3c",x"00",x"1c",x"3c"),
    56 => (x"60",x"30",x"60",x"7c"),
    57 => (x"44",x"00",x"3c",x"7c"),
    58 => (x"38",x"10",x"38",x"6c"),
    59 => (x"00",x"00",x"44",x"6c"),
    60 => (x"60",x"e0",x"bc",x"1c"),
    61 => (x"00",x"00",x"1c",x"3c"),
    62 => (x"5c",x"74",x"64",x"44"),
    63 => (x"00",x"00",x"44",x"4c"),
    64 => (x"77",x"3e",x"08",x"08"),
    65 => (x"00",x"00",x"41",x"41"),
    66 => (x"7f",x"7f",x"00",x"00"),
    67 => (x"00",x"00",x"00",x"00"),
    68 => (x"3e",x"77",x"41",x"41"),
    69 => (x"02",x"00",x"08",x"08"),
    70 => (x"02",x"03",x"01",x"01"),
    71 => (x"7f",x"00",x"01",x"02"),
    72 => (x"7f",x"7f",x"7f",x"7f"),
    73 => (x"08",x"00",x"7f",x"7f"),
    74 => (x"3e",x"1c",x"1c",x"08"),
    75 => (x"7f",x"7f",x"7f",x"3e"),
    76 => (x"1c",x"3e",x"3e",x"7f"),
    77 => (x"00",x"08",x"08",x"1c"),
    78 => (x"7c",x"7c",x"18",x"10"),
    79 => (x"00",x"00",x"10",x"18"),
    80 => (x"7c",x"7c",x"30",x"10"),
    81 => (x"10",x"00",x"10",x"30"),
    82 => (x"78",x"60",x"60",x"30"),
    83 => (x"42",x"00",x"06",x"1e"),
    84 => (x"3c",x"18",x"3c",x"66"),
    85 => (x"78",x"00",x"42",x"66"),
    86 => (x"c6",x"c2",x"6a",x"38"),
    87 => (x"60",x"00",x"38",x"6c"),
    88 => (x"00",x"60",x"00",x"00"),
    89 => (x"0e",x"00",x"60",x"00"),
    90 => (x"5d",x"5c",x"5b",x"5e"),
    91 => (x"4c",x"71",x"1e",x"0e"),
    92 => (x"bf",x"dd",x"f9",x"c2"),
    93 => (x"c0",x"4b",x"c0",x"4d"),
    94 => (x"02",x"ab",x"74",x"1e"),
    95 => (x"a6",x"c4",x"87",x"c7"),
    96 => (x"c5",x"78",x"c0",x"48"),
    97 => (x"48",x"a6",x"c4",x"87"),
    98 => (x"66",x"c4",x"78",x"c1"),
    99 => (x"ee",x"49",x"73",x"1e"),
   100 => (x"86",x"c8",x"87",x"df"),
   101 => (x"ef",x"49",x"e0",x"c0"),
   102 => (x"a5",x"c4",x"87",x"ee"),
   103 => (x"f0",x"49",x"6a",x"4a"),
   104 => (x"c6",x"f1",x"87",x"f0"),
   105 => (x"c1",x"85",x"cb",x"87"),
   106 => (x"ab",x"b7",x"c8",x"83"),
   107 => (x"87",x"c7",x"ff",x"04"),
   108 => (x"26",x"4d",x"26",x"26"),
   109 => (x"26",x"4b",x"26",x"4c"),
   110 => (x"4a",x"71",x"1e",x"4f"),
   111 => (x"5a",x"e1",x"f9",x"c2"),
   112 => (x"48",x"e1",x"f9",x"c2"),
   113 => (x"fe",x"49",x"78",x"c7"),
   114 => (x"4f",x"26",x"87",x"dd"),
   115 => (x"71",x"1e",x"73",x"1e"),
   116 => (x"aa",x"b7",x"c0",x"4a"),
   117 => (x"c2",x"87",x"d3",x"03"),
   118 => (x"05",x"bf",x"de",x"d9"),
   119 => (x"4b",x"c1",x"87",x"c4"),
   120 => (x"4b",x"c0",x"87",x"c2"),
   121 => (x"5b",x"e2",x"d9",x"c2"),
   122 => (x"d9",x"c2",x"87",x"c4"),
   123 => (x"d9",x"c2",x"5a",x"e2"),
   124 => (x"c1",x"4a",x"bf",x"de"),
   125 => (x"a2",x"c0",x"c1",x"9a"),
   126 => (x"87",x"e8",x"ec",x"49"),
   127 => (x"bf",x"c6",x"d9",x"c2"),
   128 => (x"de",x"d9",x"c2",x"48"),
   129 => (x"08",x"fc",x"b0",x"bf"),
   130 => (x"87",x"e9",x"fe",x"78"),
   131 => (x"c4",x"4a",x"71",x"1e"),
   132 => (x"49",x"72",x"1e",x"66"),
   133 => (x"26",x"87",x"f3",x"ea"),
   134 => (x"ff",x"1e",x"4f",x"26"),
   135 => (x"ff",x"c3",x"48",x"d4"),
   136 => (x"48",x"d0",x"ff",x"78"),
   137 => (x"ff",x"78",x"e1",x"c0"),
   138 => (x"78",x"c1",x"48",x"d4"),
   139 => (x"30",x"c4",x"48",x"71"),
   140 => (x"78",x"08",x"d4",x"ff"),
   141 => (x"c0",x"48",x"d0",x"ff"),
   142 => (x"4f",x"26",x"78",x"e0"),
   143 => (x"5c",x"5b",x"5e",x"0e"),
   144 => (x"86",x"f4",x"0e",x"5d"),
   145 => (x"c0",x"48",x"a6",x"c4"),
   146 => (x"bf",x"ec",x"4b",x"78"),
   147 => (x"dd",x"f9",x"c2",x"7e"),
   148 => (x"bf",x"e8",x"4d",x"bf"),
   149 => (x"de",x"d9",x"c2",x"4c"),
   150 => (x"f1",x"e3",x"49",x"bf"),
   151 => (x"49",x"f7",x"c1",x"87"),
   152 => (x"70",x"87",x"f5",x"e6"),
   153 => (x"87",x"d5",x"02",x"98"),
   154 => (x"bf",x"de",x"d9",x"c2"),
   155 => (x"87",x"de",x"e3",x"49"),
   156 => (x"f7",x"c1",x"4b",x"c1"),
   157 => (x"87",x"e0",x"e6",x"49"),
   158 => (x"eb",x"05",x"98",x"70"),
   159 => (x"02",x"9b",x"73",x"87"),
   160 => (x"c2",x"87",x"fa",x"c0"),
   161 => (x"05",x"bf",x"c6",x"d9"),
   162 => (x"a6",x"c8",x"87",x"c7"),
   163 => (x"c5",x"78",x"c1",x"48"),
   164 => (x"48",x"a6",x"c8",x"87"),
   165 => (x"d9",x"c2",x"78",x"c0"),
   166 => (x"66",x"c8",x"48",x"c6"),
   167 => (x"1e",x"fc",x"ca",x"78"),
   168 => (x"c9",x"02",x"66",x"cc"),
   169 => (x"48",x"a6",x"cc",x"87"),
   170 => (x"78",x"d9",x"d7",x"c2"),
   171 => (x"a6",x"cc",x"87",x"c7"),
   172 => (x"e4",x"d7",x"c2",x"48"),
   173 => (x"49",x"66",x"cc",x"78"),
   174 => (x"c4",x"87",x"f5",x"cc"),
   175 => (x"cb",x"4b",x"c0",x"86"),
   176 => (x"e1",x"ce",x"49",x"ee"),
   177 => (x"58",x"a6",x"cc",x"87"),
   178 => (x"cb",x"e5",x"49",x"c7"),
   179 => (x"05",x"98",x"70",x"87"),
   180 => (x"49",x"6e",x"87",x"c8"),
   181 => (x"c1",x"02",x"99",x"c1"),
   182 => (x"4b",x"c1",x"87",x"c3"),
   183 => (x"c2",x"7e",x"bf",x"ec"),
   184 => (x"49",x"bf",x"de",x"d9"),
   185 => (x"c8",x"87",x"e7",x"e1"),
   186 => (x"c5",x"ce",x"49",x"66"),
   187 => (x"02",x"98",x"70",x"87"),
   188 => (x"d9",x"c2",x"87",x"d8"),
   189 => (x"c1",x"49",x"bf",x"c2"),
   190 => (x"c6",x"d9",x"c2",x"b9"),
   191 => (x"d9",x"fc",x"71",x"59"),
   192 => (x"49",x"ee",x"cb",x"87"),
   193 => (x"cc",x"87",x"df",x"cd"),
   194 => (x"49",x"c7",x"58",x"a6"),
   195 => (x"70",x"87",x"c9",x"e4"),
   196 => (x"c5",x"ff",x"05",x"98"),
   197 => (x"c1",x"49",x"6e",x"87"),
   198 => (x"fd",x"fe",x"05",x"99"),
   199 => (x"02",x"9b",x"73",x"87"),
   200 => (x"49",x"ff",x"87",x"d0"),
   201 => (x"c1",x"87",x"e5",x"fa"),
   202 => (x"eb",x"e3",x"49",x"da"),
   203 => (x"48",x"a6",x"c4",x"87"),
   204 => (x"d9",x"c2",x"78",x"c1"),
   205 => (x"c1",x"05",x"bf",x"de"),
   206 => (x"d9",x"c2",x"87",x"e2"),
   207 => (x"c0",x"02",x"bf",x"c6"),
   208 => (x"a6",x"c4",x"87",x"f1"),
   209 => (x"c0",x"c0",x"c8",x"48"),
   210 => (x"ca",x"d9",x"c2",x"78"),
   211 => (x"bf",x"97",x"6e",x"7e"),
   212 => (x"c1",x"48",x"6e",x"49"),
   213 => (x"71",x"7e",x"70",x"80"),
   214 => (x"70",x"87",x"fd",x"e2"),
   215 => (x"c3",x"c0",x"02",x"98"),
   216 => (x"b4",x"66",x"c4",x"87"),
   217 => (x"c1",x"48",x"66",x"c4"),
   218 => (x"a6",x"c8",x"28",x"b7"),
   219 => (x"05",x"98",x"70",x"58"),
   220 => (x"c3",x"87",x"da",x"ff"),
   221 => (x"df",x"e2",x"49",x"fd"),
   222 => (x"49",x"fa",x"c3",x"87"),
   223 => (x"74",x"87",x"d9",x"e2"),
   224 => (x"99",x"ff",x"c3",x"49"),
   225 => (x"49",x"c0",x"1e",x"71"),
   226 => (x"74",x"87",x"c1",x"fa"),
   227 => (x"29",x"b7",x"c8",x"49"),
   228 => (x"49",x"c1",x"1e",x"71"),
   229 => (x"c8",x"87",x"f5",x"f9"),
   230 => (x"87",x"f8",x"c8",x"86"),
   231 => (x"ff",x"c3",x"49",x"74"),
   232 => (x"2c",x"b7",x"c8",x"99"),
   233 => (x"9c",x"74",x"b4",x"71"),
   234 => (x"87",x"e0",x"c0",x"02"),
   235 => (x"bf",x"da",x"d9",x"c2"),
   236 => (x"87",x"fe",x"ca",x"49"),
   237 => (x"c0",x"05",x"98",x"70"),
   238 => (x"4c",x"c0",x"87",x"c5"),
   239 => (x"c2",x"87",x"d3",x"c0"),
   240 => (x"e1",x"ca",x"49",x"e0"),
   241 => (x"de",x"d9",x"c2",x"87"),
   242 => (x"87",x"c6",x"c0",x"58"),
   243 => (x"48",x"da",x"d9",x"c2"),
   244 => (x"49",x"74",x"78",x"c0"),
   245 => (x"c0",x"05",x"99",x"c2"),
   246 => (x"eb",x"c3",x"87",x"ce"),
   247 => (x"87",x"f8",x"e0",x"49"),
   248 => (x"99",x"c2",x"49",x"70"),
   249 => (x"87",x"ce",x"c0",x"02"),
   250 => (x"4a",x"a5",x"d8",x"c1"),
   251 => (x"c5",x"c0",x"02",x"6a"),
   252 => (x"49",x"fb",x"4b",x"87"),
   253 => (x"49",x"74",x"0f",x"73"),
   254 => (x"c0",x"05",x"99",x"c1"),
   255 => (x"f4",x"c3",x"87",x"ce"),
   256 => (x"87",x"d4",x"e0",x"49"),
   257 => (x"99",x"c2",x"49",x"70"),
   258 => (x"87",x"cf",x"c0",x"02"),
   259 => (x"7e",x"a5",x"d8",x"c1"),
   260 => (x"c0",x"02",x"bf",x"6e"),
   261 => (x"fa",x"4b",x"87",x"c5"),
   262 => (x"74",x"0f",x"73",x"49"),
   263 => (x"05",x"99",x"c8",x"49"),
   264 => (x"c3",x"87",x"cf",x"c0"),
   265 => (x"df",x"ff",x"49",x"f5"),
   266 => (x"49",x"70",x"87",x"ee"),
   267 => (x"c0",x"02",x"99",x"c2"),
   268 => (x"f9",x"c2",x"87",x"e6"),
   269 => (x"c0",x"02",x"bf",x"e1"),
   270 => (x"c1",x"48",x"87",x"ca"),
   271 => (x"e5",x"f9",x"c2",x"88"),
   272 => (x"87",x"cf",x"c0",x"58"),
   273 => (x"7e",x"a5",x"d8",x"c1"),
   274 => (x"c0",x"02",x"bf",x"6e"),
   275 => (x"ff",x"4b",x"87",x"c5"),
   276 => (x"c4",x"0f",x"73",x"49"),
   277 => (x"78",x"c1",x"48",x"a6"),
   278 => (x"99",x"c4",x"49",x"74"),
   279 => (x"87",x"cf",x"c0",x"05"),
   280 => (x"ff",x"49",x"f2",x"c3"),
   281 => (x"70",x"87",x"f1",x"de"),
   282 => (x"02",x"99",x"c2",x"49"),
   283 => (x"c2",x"87",x"ec",x"c0"),
   284 => (x"7e",x"bf",x"e1",x"f9"),
   285 => (x"a8",x"b7",x"c7",x"48"),
   286 => (x"87",x"cb",x"c0",x"03"),
   287 => (x"80",x"c1",x"48",x"6e"),
   288 => (x"58",x"e5",x"f9",x"c2"),
   289 => (x"c1",x"87",x"cf",x"c0"),
   290 => (x"6e",x"7e",x"a5",x"d8"),
   291 => (x"c5",x"c0",x"02",x"bf"),
   292 => (x"49",x"fe",x"4b",x"87"),
   293 => (x"a6",x"c4",x"0f",x"73"),
   294 => (x"c3",x"78",x"c1",x"48"),
   295 => (x"dd",x"ff",x"49",x"fd"),
   296 => (x"49",x"70",x"87",x"f6"),
   297 => (x"c0",x"02",x"99",x"c2"),
   298 => (x"f9",x"c2",x"87",x"e5"),
   299 => (x"c0",x"02",x"bf",x"e1"),
   300 => (x"f9",x"c2",x"87",x"c9"),
   301 => (x"78",x"c0",x"48",x"e1"),
   302 => (x"c1",x"87",x"cf",x"c0"),
   303 => (x"6e",x"7e",x"a5",x"d8"),
   304 => (x"c5",x"c0",x"02",x"bf"),
   305 => (x"49",x"fd",x"4b",x"87"),
   306 => (x"a6",x"c4",x"0f",x"73"),
   307 => (x"c3",x"78",x"c1",x"48"),
   308 => (x"dd",x"ff",x"49",x"fa"),
   309 => (x"49",x"70",x"87",x"c2"),
   310 => (x"c0",x"02",x"99",x"c2"),
   311 => (x"f9",x"c2",x"87",x"e9"),
   312 => (x"c7",x"48",x"bf",x"e1"),
   313 => (x"c0",x"03",x"a8",x"b7"),
   314 => (x"f9",x"c2",x"87",x"c9"),
   315 => (x"78",x"c7",x"48",x"e1"),
   316 => (x"c1",x"87",x"cf",x"c0"),
   317 => (x"6e",x"7e",x"a5",x"d8"),
   318 => (x"c5",x"c0",x"02",x"bf"),
   319 => (x"49",x"fc",x"4b",x"87"),
   320 => (x"a6",x"c4",x"0f",x"73"),
   321 => (x"c0",x"78",x"c1",x"48"),
   322 => (x"dc",x"f9",x"c2",x"4b"),
   323 => (x"cb",x"50",x"c0",x"48"),
   324 => (x"d1",x"c5",x"49",x"ee"),
   325 => (x"58",x"a6",x"cc",x"87"),
   326 => (x"97",x"dc",x"f9",x"c2"),
   327 => (x"de",x"c1",x"05",x"bf"),
   328 => (x"c3",x"49",x"74",x"87"),
   329 => (x"c0",x"05",x"99",x"f0"),
   330 => (x"da",x"c1",x"87",x"cd"),
   331 => (x"e7",x"db",x"ff",x"49"),
   332 => (x"02",x"98",x"70",x"87"),
   333 => (x"c1",x"87",x"c8",x"c1"),
   334 => (x"4c",x"bf",x"e8",x"4b"),
   335 => (x"99",x"ff",x"c3",x"49"),
   336 => (x"71",x"2c",x"b7",x"c8"),
   337 => (x"de",x"d9",x"c2",x"b4"),
   338 => (x"d8",x"ff",x"49",x"bf"),
   339 => (x"66",x"c8",x"87",x"c0"),
   340 => (x"87",x"de",x"c4",x"49"),
   341 => (x"c0",x"02",x"98",x"70"),
   342 => (x"f9",x"c2",x"87",x"c6"),
   343 => (x"50",x"c1",x"48",x"dc"),
   344 => (x"97",x"dc",x"f9",x"c2"),
   345 => (x"d6",x"c0",x"05",x"bf"),
   346 => (x"c3",x"49",x"74",x"87"),
   347 => (x"ff",x"05",x"99",x"f0"),
   348 => (x"da",x"c1",x"87",x"c5"),
   349 => (x"df",x"da",x"ff",x"49"),
   350 => (x"05",x"98",x"70",x"87"),
   351 => (x"73",x"87",x"f8",x"fe"),
   352 => (x"dc",x"c0",x"02",x"9b"),
   353 => (x"48",x"a6",x"c8",x"87"),
   354 => (x"bf",x"e1",x"f9",x"c2"),
   355 => (x"49",x"66",x"c8",x"78"),
   356 => (x"a1",x"75",x"91",x"cb"),
   357 => (x"02",x"bf",x"6e",x"7e"),
   358 => (x"4b",x"87",x"c6",x"c0"),
   359 => (x"73",x"49",x"66",x"c8"),
   360 => (x"02",x"66",x"c4",x"0f"),
   361 => (x"c2",x"87",x"c8",x"c0"),
   362 => (x"49",x"bf",x"e1",x"f9"),
   363 => (x"c2",x"87",x"f8",x"ee"),
   364 => (x"02",x"bf",x"e2",x"d9"),
   365 => (x"49",x"87",x"dd",x"c0"),
   366 => (x"70",x"87",x"f7",x"c2"),
   367 => (x"d3",x"c0",x"02",x"98"),
   368 => (x"e1",x"f9",x"c2",x"87"),
   369 => (x"de",x"ee",x"49",x"bf"),
   370 => (x"ef",x"49",x"c0",x"87"),
   371 => (x"d9",x"c2",x"87",x"fe"),
   372 => (x"78",x"c0",x"48",x"e2"),
   373 => (x"d8",x"ef",x"8e",x"f4"),
   374 => (x"79",x"6f",x"4a",x"87"),
   375 => (x"73",x"79",x"65",x"6b"),
   376 => (x"00",x"6e",x"6f",x"20"),
   377 => (x"6b",x"79",x"6f",x"4a"),
   378 => (x"20",x"73",x"79",x"65"),
   379 => (x"00",x"66",x"66",x"6f"),
   380 => (x"5c",x"5b",x"5e",x"0e"),
   381 => (x"71",x"1e",x"0e",x"5d"),
   382 => (x"dd",x"f9",x"c2",x"4c"),
   383 => (x"cd",x"c1",x"49",x"bf"),
   384 => (x"d1",x"c1",x"4d",x"a1"),
   385 => (x"74",x"7e",x"69",x"81"),
   386 => (x"87",x"cf",x"02",x"9c"),
   387 => (x"74",x"4b",x"a5",x"c4"),
   388 => (x"dd",x"f9",x"c2",x"7b"),
   389 => (x"e0",x"ee",x"49",x"bf"),
   390 => (x"74",x"7b",x"6e",x"87"),
   391 => (x"87",x"c4",x"05",x"9c"),
   392 => (x"87",x"c2",x"4b",x"c0"),
   393 => (x"49",x"73",x"4b",x"c1"),
   394 => (x"d4",x"87",x"e1",x"ee"),
   395 => (x"87",x"c8",x"02",x"66"),
   396 => (x"87",x"f2",x"c0",x"49"),
   397 => (x"87",x"c2",x"4a",x"70"),
   398 => (x"d9",x"c2",x"4a",x"c0"),
   399 => (x"ed",x"26",x"5a",x"e6"),
   400 => (x"00",x"00",x"87",x"ef"),
   401 => (x"00",x"00",x"00",x"00"),
   402 => (x"12",x"58",x"00",x"00"),
   403 => (x"1b",x"1d",x"14",x"11"),
   404 => (x"59",x"5a",x"23",x"1c"),
   405 => (x"f2",x"f5",x"94",x"91"),
   406 => (x"00",x"00",x"f4",x"eb"),
   407 => (x"00",x"00",x"00",x"00"),
   408 => (x"00",x"00",x"00",x"00"),
   409 => (x"71",x"1e",x"00",x"00"),
   410 => (x"bf",x"c8",x"ff",x"4a"),
   411 => (x"48",x"a1",x"72",x"49"),
   412 => (x"ff",x"1e",x"4f",x"26"),
   413 => (x"fe",x"89",x"bf",x"c8"),
   414 => (x"c0",x"c0",x"c0",x"c0"),
   415 => (x"c4",x"01",x"a9",x"c0"),
   416 => (x"c2",x"4a",x"c0",x"87"),
   417 => (x"72",x"4a",x"c1",x"87"),
   418 => (x"0e",x"4f",x"26",x"48"),
   419 => (x"5d",x"5c",x"5b",x"5e"),
   420 => (x"ff",x"4b",x"71",x"0e"),
   421 => (x"66",x"d0",x"4c",x"d4"),
   422 => (x"d6",x"78",x"c0",x"48"),
   423 => (x"ef",x"d7",x"ff",x"49"),
   424 => (x"7c",x"ff",x"c3",x"87"),
   425 => (x"ff",x"c3",x"49",x"6c"),
   426 => (x"49",x"4d",x"71",x"99"),
   427 => (x"c1",x"99",x"f0",x"c3"),
   428 => (x"cb",x"05",x"a9",x"e0"),
   429 => (x"7c",x"ff",x"c3",x"87"),
   430 => (x"98",x"c3",x"48",x"6c"),
   431 => (x"78",x"08",x"66",x"d0"),
   432 => (x"6c",x"7c",x"ff",x"c3"),
   433 => (x"31",x"c8",x"49",x"4a"),
   434 => (x"6c",x"7c",x"ff",x"c3"),
   435 => (x"72",x"b2",x"71",x"4a"),
   436 => (x"c3",x"31",x"c8",x"49"),
   437 => (x"4a",x"6c",x"7c",x"ff"),
   438 => (x"49",x"72",x"b2",x"71"),
   439 => (x"ff",x"c3",x"31",x"c8"),
   440 => (x"71",x"4a",x"6c",x"7c"),
   441 => (x"48",x"d0",x"ff",x"b2"),
   442 => (x"73",x"78",x"e0",x"c0"),
   443 => (x"87",x"c2",x"02",x"9b"),
   444 => (x"48",x"75",x"7b",x"72"),
   445 => (x"4c",x"26",x"4d",x"26"),
   446 => (x"4f",x"26",x"4b",x"26"),
   447 => (x"0e",x"4f",x"26",x"1e"),
   448 => (x"0e",x"5c",x"5b",x"5e"),
   449 => (x"1e",x"76",x"86",x"f8"),
   450 => (x"fd",x"49",x"a6",x"c8"),
   451 => (x"86",x"c4",x"87",x"fd"),
   452 => (x"48",x"6e",x"4b",x"70"),
   453 => (x"c2",x"03",x"a8",x"c2"),
   454 => (x"4a",x"73",x"87",x"f0"),
   455 => (x"c1",x"9a",x"f0",x"c3"),
   456 => (x"c7",x"02",x"aa",x"d0"),
   457 => (x"aa",x"e0",x"c1",x"87"),
   458 => (x"87",x"de",x"c2",x"05"),
   459 => (x"99",x"c8",x"49",x"73"),
   460 => (x"ff",x"87",x"c3",x"02"),
   461 => (x"4c",x"73",x"87",x"c6"),
   462 => (x"ac",x"c2",x"9c",x"c3"),
   463 => (x"87",x"c2",x"c1",x"05"),
   464 => (x"c9",x"49",x"66",x"c4"),
   465 => (x"c4",x"1e",x"71",x"31"),
   466 => (x"92",x"d4",x"4a",x"66"),
   467 => (x"49",x"e5",x"f9",x"c2"),
   468 => (x"c9",x"fe",x"81",x"72"),
   469 => (x"49",x"d8",x"87",x"f1"),
   470 => (x"87",x"f4",x"d4",x"ff"),
   471 => (x"c2",x"1e",x"c0",x"c8"),
   472 => (x"fd",x"49",x"ce",x"e8"),
   473 => (x"ff",x"87",x"f7",x"e5"),
   474 => (x"e0",x"c0",x"48",x"d0"),
   475 => (x"ce",x"e8",x"c2",x"78"),
   476 => (x"4a",x"66",x"cc",x"1e"),
   477 => (x"f9",x"c2",x"92",x"d4"),
   478 => (x"81",x"72",x"49",x"e5"),
   479 => (x"87",x"f9",x"c7",x"fe"),
   480 => (x"ac",x"c1",x"86",x"cc"),
   481 => (x"87",x"c2",x"c1",x"05"),
   482 => (x"c9",x"49",x"66",x"c4"),
   483 => (x"c4",x"1e",x"71",x"31"),
   484 => (x"92",x"d4",x"4a",x"66"),
   485 => (x"49",x"e5",x"f9",x"c2"),
   486 => (x"c8",x"fe",x"81",x"72"),
   487 => (x"e8",x"c2",x"87",x"e9"),
   488 => (x"66",x"c8",x"1e",x"ce"),
   489 => (x"c2",x"92",x"d4",x"4a"),
   490 => (x"72",x"49",x"e5",x"f9"),
   491 => (x"fa",x"c5",x"fe",x"81"),
   492 => (x"ff",x"49",x"d7",x"87"),
   493 => (x"c8",x"87",x"d9",x"d3"),
   494 => (x"e8",x"c2",x"1e",x"c0"),
   495 => (x"e3",x"fd",x"49",x"ce"),
   496 => (x"86",x"cc",x"87",x"f5"),
   497 => (x"c0",x"48",x"d0",x"ff"),
   498 => (x"8e",x"f8",x"78",x"e0"),
   499 => (x"0e",x"87",x"e7",x"fc"),
   500 => (x"5d",x"5c",x"5b",x"5e"),
   501 => (x"ff",x"4a",x"71",x"0e"),
   502 => (x"66",x"d0",x"4c",x"d4"),
   503 => (x"ad",x"b7",x"c3",x"4d"),
   504 => (x"c0",x"87",x"c5",x"06"),
   505 => (x"87",x"e1",x"c1",x"48"),
   506 => (x"4b",x"75",x"1e",x"72"),
   507 => (x"f9",x"c2",x"93",x"d4"),
   508 => (x"49",x"73",x"83",x"e5"),
   509 => (x"87",x"c1",x"c0",x"fe"),
   510 => (x"4b",x"6b",x"83",x"c8"),
   511 => (x"c8",x"48",x"d0",x"ff"),
   512 => (x"7c",x"dd",x"78",x"e1"),
   513 => (x"ff",x"c3",x"48",x"73"),
   514 => (x"73",x"7c",x"70",x"98"),
   515 => (x"29",x"b7",x"c8",x"49"),
   516 => (x"ff",x"c3",x"48",x"71"),
   517 => (x"73",x"7c",x"70",x"98"),
   518 => (x"29",x"b7",x"d0",x"49"),
   519 => (x"ff",x"c3",x"48",x"71"),
   520 => (x"73",x"7c",x"70",x"98"),
   521 => (x"28",x"b7",x"d8",x"48"),
   522 => (x"7c",x"c0",x"7c",x"70"),
   523 => (x"7c",x"7c",x"7c",x"7c"),
   524 => (x"7c",x"7c",x"7c",x"7c"),
   525 => (x"ff",x"7c",x"7c",x"7c"),
   526 => (x"e0",x"c0",x"48",x"d0"),
   527 => (x"dc",x"1e",x"75",x"78"),
   528 => (x"f0",x"d1",x"ff",x"49"),
   529 => (x"73",x"86",x"c8",x"87"),
   530 => (x"87",x"e8",x"fa",x"48"),
   531 => (x"c4",x"4a",x"71",x"1e"),
   532 => (x"f9",x"c2",x"49",x"a2"),
   533 => (x"78",x"6a",x"48",x"c8"),
   534 => (x"48",x"c2",x"d9",x"c2"),
   535 => (x"d9",x"c2",x"78",x"69"),
   536 => (x"e6",x"49",x"bf",x"c2"),
   537 => (x"d1",x"ff",x"87",x"f4"),
   538 => (x"4f",x"26",x"87",x"fd"),
   539 => (x"c4",x"4a",x"71",x"1e"),
   540 => (x"f9",x"c2",x"49",x"a2"),
   541 => (x"c2",x"7a",x"bf",x"c8"),
   542 => (x"79",x"bf",x"c2",x"d9"),
   543 => (x"71",x"1e",x"4f",x"26"),
   544 => (x"c0",x"02",x"9a",x"4a"),
   545 => (x"c2",x"1e",x"87",x"ee"),
   546 => (x"fd",x"49",x"c4",x"f5"),
   547 => (x"c4",x"87",x"ea",x"fd"),
   548 => (x"02",x"98",x"70",x"86"),
   549 => (x"e8",x"c2",x"87",x"de"),
   550 => (x"f5",x"c2",x"1e",x"ce"),
   551 => (x"c2",x"fe",x"49",x"c4"),
   552 => (x"86",x"c4",x"87",x"c9"),
   553 => (x"cb",x"02",x"98",x"70"),
   554 => (x"ce",x"e8",x"c2",x"87"),
   555 => (x"87",x"dc",x"fe",x"49"),
   556 => (x"87",x"c2",x"48",x"c1"),
   557 => (x"4f",x"26",x"48",x"c0"),
   558 => (x"9a",x"4a",x"71",x"1e"),
   559 => (x"87",x"ee",x"c0",x"02"),
   560 => (x"c4",x"f5",x"c2",x"1e"),
   561 => (x"f0",x"fc",x"fd",x"49"),
   562 => (x"70",x"86",x"c4",x"87"),
   563 => (x"87",x"de",x"02",x"98"),
   564 => (x"49",x"ce",x"e8",x"c2"),
   565 => (x"c2",x"87",x"d5",x"fe"),
   566 => (x"c2",x"1e",x"ce",x"e8"),
   567 => (x"fe",x"49",x"c4",x"f5"),
   568 => (x"c4",x"87",x"d6",x"c2"),
   569 => (x"02",x"98",x"70",x"86"),
   570 => (x"48",x"c1",x"87",x"c4"),
   571 => (x"48",x"c0",x"87",x"c2"),
   572 => (x"c1",x"1e",x"4f",x"26"),
   573 => (x"c0",x"48",x"cc",x"e7"),
   574 => (x"cd",x"fa",x"c2",x"50"),
   575 => (x"87",x"cc",x"05",x"bf"),
   576 => (x"49",x"ff",x"e4",x"c2"),
   577 => (x"87",x"e1",x"d5",x"fe"),
   578 => (x"58",x"d1",x"fa",x"c2"),
   579 => (x"48",x"cc",x"e7",x"c1"),
   580 => (x"fa",x"c2",x"50",x"c2"),
   581 => (x"cc",x"05",x"bf",x"d1"),
   582 => (x"cb",x"e5",x"c2",x"87"),
   583 => (x"c8",x"d5",x"fe",x"49"),
   584 => (x"d5",x"fa",x"c2",x"87"),
   585 => (x"d5",x"fa",x"c2",x"58"),
   586 => (x"87",x"d1",x"05",x"bf"),
   587 => (x"c2",x"1e",x"f1",x"c0"),
   588 => (x"fe",x"49",x"d7",x"e5"),
   589 => (x"c4",x"87",x"c5",x"db"),
   590 => (x"d9",x"fa",x"c2",x"86"),
   591 => (x"56",x"4f",x"26",x"58"),
   592 => (x"30",x"32",x"43",x"49"),
   593 => (x"52",x"20",x"20",x"20"),
   594 => (x"4d",x"00",x"4d",x"4f"),
   595 => (x"43",x"41",x"47",x"45"),
   596 => (x"52",x"54",x"52",x"41"),
   597 => (x"4d",x"00",x"4d",x"4f"),
   598 => (x"43",x"41",x"47",x"45"),
   599 => (x"4e",x"54",x"52",x"41"),
   600 => (x"1e",x"00",x"20",x"56"),
   601 => (x"4b",x"c0",x"1e",x"73"),
   602 => (x"48",x"cd",x"fa",x"c2"),
   603 => (x"fa",x"c2",x"78",x"c0"),
   604 => (x"78",x"c0",x"48",x"d1"),
   605 => (x"48",x"d5",x"fa",x"c2"),
   606 => (x"f5",x"fd",x"78",x"c0"),
   607 => (x"d1",x"e7",x"c2",x"87"),
   608 => (x"c4",x"f5",x"c2",x"1e"),
   609 => (x"f0",x"f9",x"fd",x"49"),
   610 => (x"70",x"86",x"c4",x"87"),
   611 => (x"87",x"c9",x"02",x"98"),
   612 => (x"bf",x"c8",x"f5",x"c2"),
   613 => (x"d0",x"c2",x"fe",x"49"),
   614 => (x"87",x"d6",x"fd",x"87"),
   615 => (x"c2",x"fe",x"49",x"c0"),
   616 => (x"fa",x"c2",x"87",x"c7"),
   617 => (x"cd",x"02",x"bf",x"d1"),
   618 => (x"c8",x"f9",x"c2",x"87"),
   619 => (x"c0",x"c8",x"48",x"bf"),
   620 => (x"f9",x"c2",x"b0",x"c0"),
   621 => (x"cc",x"ff",x"58",x"cc"),
   622 => (x"fa",x"c2",x"87",x"ed"),
   623 => (x"c4",x"05",x"bf",x"cd"),
   624 => (x"dd",x"e7",x"c2",x"87"),
   625 => (x"c4",x"48",x"73",x"4b"),
   626 => (x"26",x"4d",x"26",x"87"),
   627 => (x"26",x"4b",x"26",x"4c"),
   628 => (x"41",x"48",x"43",x"4f"),
   629 => (x"20",x"30",x"32",x"4d"),
   630 => (x"20",x"20",x"20",x"20"),
   631 => (x"4d",x"4f",x"52",x"00"),
   632 => (x"69",x"61",x"66",x"20"),
   633 => (x"00",x"64",x"65",x"6c"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

