library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0d8c487",
    12 => x"86c0c84e",
    13 => x"49f0d8c4",
    14 => x"48e8fec3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087fcf1",
    19 => x"fc1e87fd",
    20 => x"ff4a7186",
    21 => x"486949c0",
    22 => x"7098c0c4",
    23 => x"0298487e",
    24 => x"797287f4",
    25 => x"268efc48",
    26 => x"1e721e4f",
    27 => x"48121e73",
    28 => x"87ca0211",
    29 => x"98dfc34b",
    30 => x"0288739b",
    31 => x"4b2687f0",
    32 => x"4f264a26",
    33 => x"721e731e",
    34 => x"048bc11e",
    35 => x"481287ca",
    36 => x"87c40211",
    37 => x"87f10288",
    38 => x"4b264a26",
    39 => x"741e4f26",
    40 => x"721e731e",
    41 => x"048bc11e",
    42 => x"481287d0",
    43 => x"87ca0211",
    44 => x"98dfc34c",
    45 => x"0288749c",
    46 => x"4a2687eb",
    47 => x"4c264b26",
    48 => x"731e4f26",
    49 => x"a9738148",
    50 => x"1287c502",
    51 => x"87f60553",
    52 => x"731e4f26",
    53 => x"a9738148",
    54 => x"f9537205",
    55 => x"1e4f2687",
    56 => x"9a721e73",
    57 => x"87e7c002",
    58 => x"4bc148c0",
    59 => x"d106a972",
    60 => x"06827287",
    61 => x"837387c9",
    62 => x"f401a972",
    63 => x"c187c387",
    64 => x"a9723ab2",
    65 => x"80738903",
    66 => x"2b2ac107",
    67 => x"2687f305",
    68 => x"1e4f264b",
    69 => x"4dc41e75",
    70 => x"04a1b771",
    71 => x"81c1b9ff",
    72 => x"7207bdc3",
    73 => x"ff04a2b7",
    74 => x"c182c1ba",
    75 => x"eefe07bd",
    76 => x"042dc187",
    77 => x"80c1b8ff",
    78 => x"ff042d07",
    79 => x"0781c1b9",
    80 => x"4f264d26",
    81 => x"711e731e",
    82 => x"4b66c84a",
    83 => x"718bc149",
    84 => x"87cf0299",
    85 => x"d4ff4812",
    86 => x"49737808",
    87 => x"99718bc1",
    88 => x"2687f105",
    89 => x"0e4f264b",
    90 => x"0e5c5b5e",
    91 => x"d4ff4a71",
    92 => x"4b66cc4c",
    93 => x"718bc149",
    94 => x"87ce0299",
    95 => x"6c7cffc3",
    96 => x"c1497352",
    97 => x"0599718b",
    98 => x"4c2687f2",
    99 => x"4f264b26",
   100 => x"ff1e731e",
   101 => x"ffc34bd4",
   102 => x"c34a6b7b",
   103 => x"496b7bff",
   104 => x"b17232c8",
   105 => x"6b7bffc3",
   106 => x"7131c84a",
   107 => x"7bffc3b2",
   108 => x"32c8496b",
   109 => x"4871b172",
   110 => x"4f264b26",
   111 => x"5c5b5e0e",
   112 => x"4d710e5d",
   113 => x"754cd4ff",
   114 => x"98ffc348",
   115 => x"fec37c70",
   116 => x"c805bfe8",
   117 => x"4866d087",
   118 => x"a6d430c9",
   119 => x"4966d058",
   120 => x"487129d8",
   121 => x"7098ffc3",
   122 => x"4966d07c",
   123 => x"487129d0",
   124 => x"7098ffc3",
   125 => x"4966d07c",
   126 => x"487129c8",
   127 => x"7098ffc3",
   128 => x"4866d07c",
   129 => x"7098ffc3",
   130 => x"d049757c",
   131 => x"c3487129",
   132 => x"7c7098ff",
   133 => x"f0c94b6c",
   134 => x"ffc34aff",
   135 => x"87cf05ab",
   136 => x"6c7c7149",
   137 => x"028ac14b",
   138 => x"ab7187c5",
   139 => x"7387f202",
   140 => x"264d2648",
   141 => x"264b264c",
   142 => x"49c01e4f",
   143 => x"c348d4ff",
   144 => x"81c178ff",
   145 => x"a9b7c8c3",
   146 => x"2687f104",
   147 => x"5b5e0e4f",
   148 => x"c00e5d5c",
   149 => x"f7c1f0ff",
   150 => x"c0c0c14d",
   151 => x"4bc0c0c0",
   152 => x"c487d6ff",
   153 => x"c04cdff8",
   154 => x"fd49751e",
   155 => x"86c487ce",
   156 => x"c005a8c1",
   157 => x"d4ff87e5",
   158 => x"78ffc348",
   159 => x"e1c01e73",
   160 => x"49e9c1f0",
   161 => x"c487f5fc",
   162 => x"05987086",
   163 => x"d4ff87ca",
   164 => x"78ffc348",
   165 => x"87cb48c1",
   166 => x"c187defe",
   167 => x"c6ff058c",
   168 => x"2648c087",
   169 => x"264c264d",
   170 => x"0e4f264b",
   171 => x"0e5c5b5e",
   172 => x"c1f0ffc0",
   173 => x"d4ff4cc1",
   174 => x"78ffc348",
   175 => x"1ec04bd3",
   176 => x"f7fb4974",
   177 => x"7086c487",
   178 => x"87ca0598",
   179 => x"c348d4ff",
   180 => x"48c178ff",
   181 => x"e0fd87ca",
   182 => x"058bc187",
   183 => x"48c087e0",
   184 => x"4b264c26",
   185 => x"5e0e4f26",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"c4fd4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"fbfa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087e0fe",
   195 => x"87e2c148",
   196 => x"7087fdf9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fe87c802",
   200 => x"48c087c9",
   201 => x"7587cbc1",
   202 => x"4cf1c07b",
   203 => x"7087defc",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87fcf949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"d548c187",
   215 => x"d148c087",
   216 => x"05acc287",
   217 => x"48c087c4",
   218 => x"8cc187c8",
   219 => x"87fcfe05",
   220 => x"4d2648c0",
   221 => x"4b264c26",
   222 => x"5e0e4f26",
   223 => x"0e5d5c5b",
   224 => x"c04dd0ff",
   225 => x"c0c1d0e5",
   226 => x"e8fec34c",
   227 => x"c778c148",
   228 => x"fa7dc24b",
   229 => x"7dc387e3",
   230 => x"49741ec0",
   231 => x"c487ddf8",
   232 => x"05a8c186",
   233 => x"c24b87c1",
   234 => x"87c505ab",
   235 => x"f6c048c0",
   236 => x"058bc187",
   237 => x"fc87daff",
   238 => x"fec387ec",
   239 => x"987058ec",
   240 => x"c187cd05",
   241 => x"f0ffc01e",
   242 => x"f749d0c1",
   243 => x"86c487ee",
   244 => x"c348d4ff",
   245 => x"e8c478ff",
   246 => x"f0fec387",
   247 => x"ff7dc258",
   248 => x"ffc348d4",
   249 => x"2648c178",
   250 => x"264c264d",
   251 => x"0e4f264b",
   252 => x"5d5c5b5e",
   253 => x"c34d710e",
   254 => x"d4ff4cff",
   255 => x"ff7b744b",
   256 => x"c3c448d0",
   257 => x"757b7478",
   258 => x"f0ffc01e",
   259 => x"f649d8c1",
   260 => x"86c487ea",
   261 => x"c5029870",
   262 => x"c048c187",
   263 => x"7b7487ee",
   264 => x"c87bfec3",
   265 => x"66d41ec0",
   266 => x"87d8f449",
   267 => x"7b7486c4",
   268 => x"7b747b74",
   269 => x"4ae0dad8",
   270 => x"056b7b74",
   271 => x"8ac187c5",
   272 => x"7487f505",
   273 => x"48d0ff7b",
   274 => x"48c078c2",
   275 => x"4c264d26",
   276 => x"4f264b26",
   277 => x"5c5b5e0e",
   278 => x"86fc0e5d",
   279 => x"d4ff4b71",
   280 => x"c57ec04c",
   281 => x"4adfcdee",
   282 => x"6c7cffc3",
   283 => x"a8fec348",
   284 => x"87f8c005",
   285 => x"9b734d74",
   286 => x"d487cc02",
   287 => x"49731e66",
   288 => x"c487e4f3",
   289 => x"ff87d486",
   290 => x"d1c448d0",
   291 => x"4a66d478",
   292 => x"c17dffc3",
   293 => x"87f8058a",
   294 => x"c35aa6d8",
   295 => x"737c7cff",
   296 => x"87c5059b",
   297 => x"d048d0ff",
   298 => x"7e4ac178",
   299 => x"fe058ac1",
   300 => x"486e87f6",
   301 => x"4d268efc",
   302 => x"4b264c26",
   303 => x"731e4f26",
   304 => x"c04a711e",
   305 => x"48d4ff4b",
   306 => x"ff78ffc3",
   307 => x"c3c448d0",
   308 => x"48d4ff78",
   309 => x"7278ffc3",
   310 => x"f0ffc01e",
   311 => x"f349d1c1",
   312 => x"86c487da",
   313 => x"d2059870",
   314 => x"1ec0c887",
   315 => x"fd4966cc",
   316 => x"86c487e2",
   317 => x"d0ff4b70",
   318 => x"7378c248",
   319 => x"264b2648",
   320 => x"5b5e0e4f",
   321 => x"c00e5d5c",
   322 => x"f0ffc01e",
   323 => x"f249c9c1",
   324 => x"1ed287ea",
   325 => x"49f0fec3",
   326 => x"c887f9fc",
   327 => x"c14cc086",
   328 => x"acb7d284",
   329 => x"c387f804",
   330 => x"bf97f0fe",
   331 => x"99c0c349",
   332 => x"05a9c0c1",
   333 => x"c387e7c0",
   334 => x"bf97f7fe",
   335 => x"c331d049",
   336 => x"bf97f8fe",
   337 => x"7232c84a",
   338 => x"f9fec3b1",
   339 => x"b14abf97",
   340 => x"ffcf4c71",
   341 => x"c19cffff",
   342 => x"c134ca84",
   343 => x"fec387e7",
   344 => x"49bf97f9",
   345 => x"99c631c1",
   346 => x"97fafec3",
   347 => x"b7c74abf",
   348 => x"c3b1722a",
   349 => x"bf97f5fe",
   350 => x"9dcf4d4a",
   351 => x"97f6fec3",
   352 => x"9ac34abf",
   353 => x"fec332ca",
   354 => x"4bbf97f7",
   355 => x"b27333c2",
   356 => x"97f8fec3",
   357 => x"c0c34bbf",
   358 => x"2bb7c69b",
   359 => x"81c2b273",
   360 => x"307148c1",
   361 => x"48c14970",
   362 => x"4d703075",
   363 => x"84c14c72",
   364 => x"c0c89471",
   365 => x"cc06adb7",
   366 => x"b734c187",
   367 => x"b7c0c82d",
   368 => x"f4ff01ad",
   369 => x"26487487",
   370 => x"264c264d",
   371 => x"0e4f264b",
   372 => x"5d5c5b5e",
   373 => x"c486f80e",
   374 => x"c048d8c7",
   375 => x"d0ffc378",
   376 => x"fb49c01e",
   377 => x"86c487d8",
   378 => x"c5059870",
   379 => x"c948c087",
   380 => x"4dc087c0",
   381 => x"c2c17ec1",
   382 => x"c449bfd0",
   383 => x"714ac6c0",
   384 => x"ffe94bc8",
   385 => x"05987087",
   386 => x"7ec087c2",
   387 => x"bfccc2c1",
   388 => x"e2c0c449",
   389 => x"4bc8714a",
   390 => x"7087e9e9",
   391 => x"87c20598",
   392 => x"026e7ec0",
   393 => x"c487fdc0",
   394 => x"4dbfd6c6",
   395 => x"9fcec7c4",
   396 => x"c5487ebf",
   397 => x"05a8ead6",
   398 => x"c6c487c7",
   399 => x"ce4dbfd6",
   400 => x"ca486e87",
   401 => x"02a8d5e9",
   402 => x"48c087c5",
   403 => x"c387e3c7",
   404 => x"751ed0ff",
   405 => x"87e6f949",
   406 => x"987086c4",
   407 => x"c087c505",
   408 => x"87cec748",
   409 => x"bfccc2c1",
   410 => x"e2c0c449",
   411 => x"4bc8714a",
   412 => x"7087d1e8",
   413 => x"87c80598",
   414 => x"48d8c7c4",
   415 => x"87da78c1",
   416 => x"bfd0c2c1",
   417 => x"c6c0c449",
   418 => x"4bc8714a",
   419 => x"7087f5e7",
   420 => x"c5c00298",
   421 => x"c648c087",
   422 => x"c7c487d8",
   423 => x"49bf97ce",
   424 => x"05a9d5c1",
   425 => x"c487cdc0",
   426 => x"bf97cfc7",
   427 => x"a9eac249",
   428 => x"87c5c002",
   429 => x"f9c548c0",
   430 => x"d0ffc387",
   431 => x"487ebf97",
   432 => x"02a8e9c3",
   433 => x"6e87cec0",
   434 => x"a8ebc348",
   435 => x"87c5c002",
   436 => x"ddc548c0",
   437 => x"dbffc387",
   438 => x"9949bf97",
   439 => x"87ccc005",
   440 => x"97dcffc3",
   441 => x"a9c249bf",
   442 => x"87c5c002",
   443 => x"c1c548c0",
   444 => x"ddffc387",
   445 => x"c448bf97",
   446 => x"7058d4c7",
   447 => x"88c1484c",
   448 => x"58d8c7c4",
   449 => x"97deffc3",
   450 => x"817549bf",
   451 => x"97dfffc3",
   452 => x"32c84abf",
   453 => x"c47ea172",
   454 => x"6e48e8cb",
   455 => x"e0ffc378",
   456 => x"c848bf97",
   457 => x"c7c458a6",
   458 => x"c202bfd8",
   459 => x"c2c187cf",
   460 => x"c449bfcc",
   461 => x"714ae2c0",
   462 => x"c7e54bc8",
   463 => x"02987087",
   464 => x"c087c5c0",
   465 => x"87eac348",
   466 => x"bfd0c7c4",
   467 => x"fccbc44c",
   468 => x"f5ffc35c",
   469 => x"c849bf97",
   470 => x"f4ffc331",
   471 => x"a14abf97",
   472 => x"f6ffc349",
   473 => x"d04abf97",
   474 => x"49a17232",
   475 => x"97f7ffc3",
   476 => x"32d84abf",
   477 => x"c449a172",
   478 => x"cbc49166",
   479 => x"c481bfe8",
   480 => x"c359f0cb",
   481 => x"bf97fdff",
   482 => x"c332c84a",
   483 => x"bf97fcff",
   484 => x"c34aa24b",
   485 => x"bf97feff",
   486 => x"7333d04b",
   487 => x"ffc34aa2",
   488 => x"4bbf97ff",
   489 => x"33d89bcf",
   490 => x"c44aa273",
   491 => x"c25af4cb",
   492 => x"c492748a",
   493 => x"7248f4cb",
   494 => x"c1c178a1",
   495 => x"e2ffc387",
   496 => x"c849bf97",
   497 => x"e1ffc331",
   498 => x"a14abf97",
   499 => x"c731c549",
   500 => x"29c981ff",
   501 => x"59fccbc4",
   502 => x"97e7ffc3",
   503 => x"32c84abf",
   504 => x"97e6ffc3",
   505 => x"4aa24bbf",
   506 => x"6e9266c4",
   507 => x"f8cbc482",
   508 => x"f0cbc45a",
   509 => x"c478c048",
   510 => x"7248eccb",
   511 => x"cbc478a1",
   512 => x"cbc448fc",
   513 => x"c478bff0",
   514 => x"c448c0cc",
   515 => x"78bff4cb",
   516 => x"bfd8c7c4",
   517 => x"87c9c002",
   518 => x"30c44874",
   519 => x"c9c07e70",
   520 => x"f8cbc487",
   521 => x"30c448bf",
   522 => x"c7c47e70",
   523 => x"786e48dc",
   524 => x"8ef848c1",
   525 => x"4c264d26",
   526 => x"4f264b26",
   527 => x"5c5b5e0e",
   528 => x"4a710e5d",
   529 => x"bfd8c7c4",
   530 => x"7287cb02",
   531 => x"722bc74b",
   532 => x"9dffc14d",
   533 => x"4b7287c9",
   534 => x"4d722bc8",
   535 => x"c49dffc3",
   536 => x"83bfe8cb",
   537 => x"bfc8c2c1",
   538 => x"87d902ab",
   539 => x"5bccc2c1",
   540 => x"1ed0ffc3",
   541 => x"c5f14973",
   542 => x"7086c487",
   543 => x"87c50598",
   544 => x"e6c048c0",
   545 => x"d8c7c487",
   546 => x"87d202bf",
   547 => x"91c44975",
   548 => x"81d0ffc3",
   549 => x"ffcf4c69",
   550 => x"9cffffff",
   551 => x"497587cb",
   552 => x"ffc391c2",
   553 => x"699f81d0",
   554 => x"2648744c",
   555 => x"264c264d",
   556 => x"0e4f264b",
   557 => x"5d5c5b5e",
   558 => x"cc86f00e",
   559 => x"66c859a6",
   560 => x"c087c505",
   561 => x"87c4c448",
   562 => x"c84866c8",
   563 => x"487e7080",
   564 => x"e0c078c0",
   565 => x"87c80266",
   566 => x"9766e0c0",
   567 => x"87c505bf",
   568 => x"e7c348c0",
   569 => x"c11ec087",
   570 => x"c2d14949",
   571 => x"7086c487",
   572 => x"c0029c4c",
   573 => x"c7c487fe",
   574 => x"e0c04ae0",
   575 => x"ddff4966",
   576 => x"987087e7",
   577 => x"87ecc002",
   578 => x"e0c04a74",
   579 => x"4bcb4966",
   580 => x"87cadeff",
   581 => x"db029870",
   582 => x"741ec087",
   583 => x"87c4029c",
   584 => x"87c24dc0",
   585 => x"49754dc1",
   586 => x"c487c4d0",
   587 => x"9c4c7086",
   588 => x"87c2ff05",
   589 => x"c2029c74",
   590 => x"a4dc87d0",
   591 => x"69486e49",
   592 => x"49a4da78",
   593 => x"c44866c8",
   594 => x"58a6c880",
   595 => x"c448699f",
   596 => x"c4780866",
   597 => x"02bfd8c7",
   598 => x"a4d487d2",
   599 => x"49699f49",
   600 => x"99ffffc0",
   601 => x"30d04871",
   602 => x"87c558a6",
   603 => x"c048a6cc",
   604 => x"4866cc78",
   605 => x"80bf66c4",
   606 => x"780866c4",
   607 => x"c04866c8",
   608 => x"4966c878",
   609 => x"66c481cc",
   610 => x"66c879bf",
   611 => x"c081d049",
   612 => x"66c44d79",
   613 => x"4a66c84c",
   614 => x"497582d4",
   615 => x"a17291c8",
   616 => x"6c41c049",
   617 => x"c685c179",
   618 => x"ff04adb7",
   619 => x"bf6e87e7",
   620 => x"722ac94a",
   621 => x"4af0c049",
   622 => x"87e3dcff",
   623 => x"66c84a70",
   624 => x"81c4c149",
   625 => x"48c17972",
   626 => x"48c087c2",
   627 => x"4d268ef0",
   628 => x"4b264c26",
   629 => x"5e0e4f26",
   630 => x"0e5d5c5b",
   631 => x"66d04c71",
   632 => x"029c744d",
   633 => x"c887c2c1",
   634 => x"026949a4",
   635 => x"6c87fac0",
   636 => x"b9758549",
   637 => x"bfd4c7c4",
   638 => x"72baff4a",
   639 => x"02997199",
   640 => x"c487e4c0",
   641 => x"496b4ba4",
   642 => x"7087f1f8",
   643 => x"d0c7c47b",
   644 => x"816c49bf",
   645 => x"b9757c71",
   646 => x"bfd4c7c4",
   647 => x"72baff4a",
   648 => x"05997199",
   649 => x"7587dcff",
   650 => x"264d267c",
   651 => x"264b264c",
   652 => x"1e731e4f",
   653 => x"029b4b71",
   654 => x"a3c887c7",
   655 => x"c5056949",
   656 => x"c048c087",
   657 => x"cbc487f6",
   658 => x"c449bfec",
   659 => x"4a6a4aa3",
   660 => x"c7c48ac2",
   661 => x"7292bfd0",
   662 => x"c7c449a1",
   663 => x"6b4abfd4",
   664 => x"49a1729a",
   665 => x"59ccc2c1",
   666 => x"711e66c8",
   667 => x"c487cfe9",
   668 => x"05987086",
   669 => x"48c087c4",
   670 => x"48c187c2",
   671 => x"4f264b26",
   672 => x"711e731e",
   673 => x"c7029b4b",
   674 => x"49a3c887",
   675 => x"87c50569",
   676 => x"f6c048c0",
   677 => x"eccbc487",
   678 => x"a3c449bf",
   679 => x"c24a6a4a",
   680 => x"d0c7c48a",
   681 => x"a17292bf",
   682 => x"d4c7c449",
   683 => x"9a6b4abf",
   684 => x"c149a172",
   685 => x"c859ccc2",
   686 => x"e4711e66",
   687 => x"86c487f1",
   688 => x"c4059870",
   689 => x"c248c087",
   690 => x"2648c187",
   691 => x"0e4f264b",
   692 => x"5d5c5b5e",
   693 => x"7186f80e",
   694 => x"48a6c47e",
   695 => x"ffc178ff",
   696 => x"ffffffff",
   697 => x"6e4bc04d",
   698 => x"7382d44a",
   699 => x"7291c849",
   700 => x"66d849a1",
   701 => x"c08c694c",
   702 => x"cb04acb7",
   703 => x"acb77587",
   704 => x"c887c503",
   705 => x"4d745ba6",
   706 => x"b7c683c1",
   707 => x"d6ff04ab",
   708 => x"4866c487",
   709 => x"4d268ef8",
   710 => x"4b264c26",
   711 => x"5e0e4f26",
   712 => x"0e5d5c5b",
   713 => x"7e7186f0",
   714 => x"c148a6c4",
   715 => x"ffffffff",
   716 => x"80c478ff",
   717 => x"4dc078ff",
   718 => x"4b6e4cc0",
   719 => x"4a7483d4",
   720 => x"a27392c8",
   721 => x"c849754a",
   722 => x"49a17391",
   723 => x"8869486a",
   724 => x"a6d04970",
   725 => x"02ad7459",
   726 => x"66cc87d2",
   727 => x"a866c448",
   728 => x"cc87c903",
   729 => x"a6c45ca6",
   730 => x"7866cc48",
   731 => x"b7c684c1",
   732 => x"c5ff04ac",
   733 => x"c685c187",
   734 => x"fe04adb7",
   735 => x"66c887fa",
   736 => x"268ef048",
   737 => x"264c264d",
   738 => x"0e4f264b",
   739 => x"5d5c5b5e",
   740 => x"7186ec0e",
   741 => x"66e4c04b",
   742 => x"c828c948",
   743 => x"c7c458a6",
   744 => x"ff4abfd4",
   745 => x"c44872ba",
   746 => x"a6cc9866",
   747 => x"029b7358",
   748 => x"c887c1c3",
   749 => x"026949a3",
   750 => x"7287f9c2",
   751 => x"d4986b48",
   752 => x"a3c458a6",
   753 => x"c87e6c4c",
   754 => x"66d04866",
   755 => x"87c605a8",
   756 => x"c27b66c4",
   757 => x"66c887cc",
   758 => x"fb49731e",
   759 => x"86c487f1",
   760 => x"b7c04d70",
   761 => x"87d004ad",
   762 => x"754aa3d4",
   763 => x"7291c849",
   764 => x"7b2149a1",
   765 => x"87c77c69",
   766 => x"a3cc7bc0",
   767 => x"c47c6949",
   768 => x"886b4866",
   769 => x"d058a6c8",
   770 => x"49731e66",
   771 => x"c487c0fb",
   772 => x"c14d7086",
   773 => x"c849a3c4",
   774 => x"786948a6",
   775 => x"c84866d0",
   776 => x"c006a866",
   777 => x"b7c087f2",
   778 => x"ebc004ad",
   779 => x"48a6cc87",
   780 => x"7578a3d4",
   781 => x"cc91c849",
   782 => x"66d08166",
   783 => x"70886948",
   784 => x"a966c849",
   785 => x"7387d106",
   786 => x"87d2fb49",
   787 => x"91c84970",
   788 => x"d08166cc",
   789 => x"796e4166",
   790 => x"731e66c4",
   791 => x"87f6f549",
   792 => x"ffc386c4",
   793 => x"49731ed0",
   794 => x"c487c6f7",
   795 => x"49a3d086",
   796 => x"7966e4c0",
   797 => x"4d268eec",
   798 => x"4b264c26",
   799 => x"731e4f26",
   800 => x"9b4b711e",
   801 => x"87e4c002",
   802 => x"5bc0ccc4",
   803 => x"8ac24a73",
   804 => x"bfd0c7c4",
   805 => x"cbc49249",
   806 => x"7248bfec",
   807 => x"c4ccc480",
   808 => x"c4487158",
   809 => x"e0c7c430",
   810 => x"87edc058",
   811 => x"48fccbc4",
   812 => x"bff0cbc4",
   813 => x"c0ccc478",
   814 => x"f4cbc448",
   815 => x"c7c478bf",
   816 => x"c902bfd8",
   817 => x"d0c7c487",
   818 => x"31c449bf",
   819 => x"cbc487c7",
   820 => x"c449bff8",
   821 => x"e0c7c431",
   822 => x"264b2659",
   823 => x"cbc41e4f",
   824 => x"c449bffc",
   825 => x"a9bff0cb",
   826 => x"c087c405",
   827 => x"7187c24a",
   828 => x"2648724a",
   829 => x"5b5e0e4f",
   830 => x"4a710e5c",
   831 => x"9a724bc0",
   832 => x"87e0c002",
   833 => x"9f49a2da",
   834 => x"c7c44b69",
   835 => x"cf02bfd8",
   836 => x"49a2d487",
   837 => x"4c49699f",
   838 => x"9cffffc0",
   839 => x"87c234d0",
   840 => x"b3744cc0",
   841 => x"d5fd4973",
   842 => x"264c2687",
   843 => x"0e4f264b",
   844 => x"5d5c5b5e",
   845 => x"c886f00e",
   846 => x"ffcf59a6",
   847 => x"4cf8ffff",
   848 => x"66c47ec0",
   849 => x"c387d802",
   850 => x"c048ccff",
   851 => x"c4ffc378",
   852 => x"c0ccc448",
   853 => x"ffc378bf",
   854 => x"cbc448c8",
   855 => x"c478bffc",
   856 => x"c048edc7",
   857 => x"dcc7c450",
   858 => x"ffc349bf",
   859 => x"714abfcc",
   860 => x"ccc403aa",
   861 => x"cf497287",
   862 => x"eac00599",
   863 => x"c8c2c187",
   864 => x"c4ffc348",
   865 => x"ffc378bf",
   866 => x"ffc31ed0",
   867 => x"c349bfc4",
   868 => x"c148c4ff",
   869 => x"ff7178a1",
   870 => x"c487e3dc",
   871 => x"e4fcc086",
   872 => x"d0ffc348",
   873 => x"c087cc78",
   874 => x"48bfe4fc",
   875 => x"c080e0c0",
   876 => x"c358e8fc",
   877 => x"48bfccff",
   878 => x"ffc380c1",
   879 => x"242758d0",
   880 => x"bf00000f",
   881 => x"9d4dbf97",
   882 => x"87e5c202",
   883 => x"02ade5c3",
   884 => x"c087dec2",
   885 => x"4bbfe4fc",
   886 => x"1149a3cb",
   887 => x"05accf4c",
   888 => x"7587d2c1",
   889 => x"c199df49",
   890 => x"c491cd89",
   891 => x"c181e0c7",
   892 => x"51124aa3",
   893 => x"124aa3c3",
   894 => x"4aa3c551",
   895 => x"a3c75112",
   896 => x"c951124a",
   897 => x"51124aa3",
   898 => x"124aa3ce",
   899 => x"4aa3d051",
   900 => x"a3d25112",
   901 => x"d451124a",
   902 => x"51124aa3",
   903 => x"124aa3d6",
   904 => x"4aa3d851",
   905 => x"a3dc5112",
   906 => x"de51124a",
   907 => x"51124aa3",
   908 => x"fcc07ec1",
   909 => x"c8497487",
   910 => x"edc00599",
   911 => x"d0497487",
   912 => x"87d30599",
   913 => x"0266e0c0",
   914 => x"7387ccc0",
   915 => x"66e0c049",
   916 => x"0298700f",
   917 => x"6e87d3c0",
   918 => x"87c6c005",
   919 => x"48e0c7c4",
   920 => x"fcc050c0",
   921 => x"c248bfe4",
   922 => x"c7c487e9",
   923 => x"50c048ed",
   924 => x"dcc7c47e",
   925 => x"ffc349bf",
   926 => x"714abfcc",
   927 => x"f4fb04aa",
   928 => x"ffffcf87",
   929 => x"c44cf8ff",
   930 => x"05bfc0cc",
   931 => x"c487c8c0",
   932 => x"02bfd8c7",
   933 => x"c387fac1",
   934 => x"49bfc8ff",
   935 => x"c387dde6",
   936 => x"c458ccff",
   937 => x"ffc348a6",
   938 => x"c478bfc8",
   939 => x"02bfd8c7",
   940 => x"c487dbc0",
   941 => x"99744966",
   942 => x"c002a974",
   943 => x"a6c887c8",
   944 => x"c078c048",
   945 => x"a6c887e7",
   946 => x"c078c148",
   947 => x"66c487df",
   948 => x"f8ffcf49",
   949 => x"c002a999",
   950 => x"a6cc87c8",
   951 => x"c078c048",
   952 => x"a6cc87c5",
   953 => x"c878c148",
   954 => x"66cc48a6",
   955 => x"0566c878",
   956 => x"c487dec0",
   957 => x"89c24966",
   958 => x"bfd0c7c4",
   959 => x"eccbc491",
   960 => x"807148bf",
   961 => x"58c8ffc3",
   962 => x"48ccffc3",
   963 => x"d4f978c0",
   964 => x"cf48c087",
   965 => x"f8ffffff",
   966 => x"268ef04c",
   967 => x"264c264d",
   968 => x"004f264b",
   969 => x"00000000",
   970 => x"5c5b5e0e",
   971 => x"86fc0e5d",
   972 => x"496e7e71",
   973 => x"c087c7f5",
   974 => x"4949c11e",
   975 => x"c487f0f7",
   976 => x"9a4a7086",
   977 => x"87c6c102",
   978 => x"9f49a2da",
   979 => x"c7c44b69",
   980 => x"cf02bfd8",
   981 => x"49a2d487",
   982 => x"4c49699f",
   983 => x"9cffffc0",
   984 => x"87c234d0",
   985 => x"a3744cc0",
   986 => x"ab66d44b",
   987 => x"c187c405",
   988 => x"c087dd48",
   989 => x"029a721e",
   990 => x"4dc087c4",
   991 => x"4dc187c2",
   992 => x"eaf64975",
   993 => x"7086c487",
   994 => x"fe059a4a",
   995 => x"48c087fa",
   996 => x"4d268efc",
   997 => x"4b264c26",
   998 => x"5e0e4f26",
   999 => x"0e5d5c5b",
  1000 => x"a6c886f4",
  1001 => x"0266c459",
  1002 => x"c44887c9",
  1003 => x"a8bff0cb",
  1004 => x"c187c505",
  1005 => x"87f7c248",
  1006 => x"c24966c4",
  1007 => x"d0c7c489",
  1008 => x"cbc491bf",
  1009 => x"c381bfec",
  1010 => x"711ed0ff",
  1011 => x"87eed3ff",
  1012 => x"987086c4",
  1013 => x"c087c505",
  1014 => x"87d3c248",
  1015 => x"4cd0ffc3",
  1016 => x"6c977ec0",
  1017 => x"58a6cc48",
  1018 => x"c1029870",
  1019 => x"c34887ef",
  1020 => x"c102a8e5",
  1021 => x"a4cb87e7",
  1022 => x"49699749",
  1023 => x"c10299d0",
  1024 => x"4a7487db",
  1025 => x"49fcc1c1",
  1026 => x"c1ff4bc8",
  1027 => x"987087f6",
  1028 => x"87c9c105",
  1029 => x"c47ea4da",
  1030 => x"02bfd8c7",
  1031 => x"a4d487cf",
  1032 => x"49699f49",
  1033 => x"ffffc04d",
  1034 => x"c235d09d",
  1035 => x"6e4dc087",
  1036 => x"7549bf9f",
  1037 => x"59a6cc81",
  1038 => x"fd4966c8",
  1039 => x"987087dc",
  1040 => x"c487d402",
  1041 => x"66cc1e66",
  1042 => x"87dcfb49",
  1043 => x"987086c4",
  1044 => x"c187c402",
  1045 => x"c087c27e",
  1046 => x"d2486e7e",
  1047 => x"84e0c087",
  1048 => x"80c1486e",
  1049 => x"d0487e70",
  1050 => x"f5fd04a8",
  1051 => x"f448c087",
  1052 => x"264d268e",
  1053 => x"264b264c",
  1054 => x"0000004f",
  1055 => x"20202e2e",
  1056 => x"20202020",
  1057 => x"00202020",
  1058 => x"ffffffff",
  1059 => x"00001094",
  1060 => x"000010a0",
  1061 => x"33544146",
  1062 => x"20202032",
  1063 => x"00000000",
  1064 => x"31544146",
  1065 => x"20202036",
  1066 => x"d0ff1e00",
  1067 => x"78e0c048",
  1068 => x"c21e4f26",
  1069 => x"7087d9d2",
  1070 => x"c6029949",
  1071 => x"a9fbc087",
  1072 => x"7187f005",
  1073 => x"0e4f2648",
  1074 => x"0e5c5b5e",
  1075 => x"4cc04b71",
  1076 => x"87fcd1c2",
  1077 => x"02994970",
  1078 => x"c087fac0",
  1079 => x"c002a9ec",
  1080 => x"fbc087f3",
  1081 => x"ecc002a9",
  1082 => x"b766cc87",
  1083 => x"87c703ac",
  1084 => x"c20266d0",
  1085 => x"71537187",
  1086 => x"87c20299",
  1087 => x"d1c284c1",
  1088 => x"497087ce",
  1089 => x"87cd0299",
  1090 => x"02a9ecc0",
  1091 => x"fbc087c7",
  1092 => x"d4ff05a9",
  1093 => x"0266d087",
  1094 => x"97c087c3",
  1095 => x"a9ecc07b",
  1096 => x"7487c405",
  1097 => x"7487c54a",
  1098 => x"8a0ac04a",
  1099 => x"4c264872",
  1100 => x"4f264b26",
  1101 => x"d7d0c21e",
  1102 => x"4a497087",
  1103 => x"04aaf0c0",
  1104 => x"f9c087c9",
  1105 => x"87c301aa",
  1106 => x"c18af0c0",
  1107 => x"c904aac1",
  1108 => x"aadac187",
  1109 => x"c087c301",
  1110 => x"48728af7",
  1111 => x"5e0e4f26",
  1112 => x"0e5d5c5b",
  1113 => x"4c7186f8",
  1114 => x"d0c27ec0",
  1115 => x"4bc087c5",
  1116 => x"97c4c8c1",
  1117 => x"a9c049bf",
  1118 => x"fc87cf04",
  1119 => x"83c187f4",
  1120 => x"97c4c8c1",
  1121 => x"06ab49bf",
  1122 => x"c8c187f1",
  1123 => x"02bf97c4",
  1124 => x"cec287d0",
  1125 => x"497087fa",
  1126 => x"87c60299",
  1127 => x"05a9ecc0",
  1128 => x"4bc087f0",
  1129 => x"87e8cec2",
  1130 => x"cec24d70",
  1131 => x"a6c887e2",
  1132 => x"dbcec258",
  1133 => x"c14a7087",
  1134 => x"49a4c883",
  1135 => x"ad496997",
  1136 => x"c987da05",
  1137 => x"699749a4",
  1138 => x"a966c449",
  1139 => x"ca87ce05",
  1140 => x"699749a4",
  1141 => x"c405aa49",
  1142 => x"d07ec187",
  1143 => x"adecc087",
  1144 => x"c087c602",
  1145 => x"c405adfb",
  1146 => x"c14bc087",
  1147 => x"fe026e7e",
  1148 => x"f4fa87f2",
  1149 => x"f8487387",
  1150 => x"264d268e",
  1151 => x"264b264c",
  1152 => x"0000004f",
  1153 => x"5b5e0e00",
  1154 => x"f40e5d5c",
  1155 => x"ff7e7186",
  1156 => x"1e6e4bd4",
  1157 => x"49ccccc4",
  1158 => x"87d7daff",
  1159 => x"987086c4",
  1160 => x"87f7c402",
  1161 => x"c148a6c4",
  1162 => x"78bfe8f3",
  1163 => x"edfc496e",
  1164 => x"58a6cc87",
  1165 => x"c5059870",
  1166 => x"48a6c887",
  1167 => x"d0ff78c1",
  1168 => x"c178c548",
  1169 => x"66c87bd5",
  1170 => x"c689c149",
  1171 => x"e0f3c131",
  1172 => x"484abf97",
  1173 => x"7b70b071",
  1174 => x"c448d0ff",
  1175 => x"c4ccc478",
  1176 => x"d049bf97",
  1177 => x"87d70299",
  1178 => x"d6c178c5",
  1179 => x"c34ac07b",
  1180 => x"82c17bff",
  1181 => x"04aae0c0",
  1182 => x"d0ff87f5",
  1183 => x"c378c448",
  1184 => x"d0ff7bff",
  1185 => x"c178c548",
  1186 => x"7bc17bd3",
  1187 => x"7e7378c4",
  1188 => x"c04866c4",
  1189 => x"c206a8b7",
  1190 => x"ccc487ee",
  1191 => x"c44cbfd4",
  1192 => x"88744866",
  1193 => x"7458a6c8",
  1194 => x"f7c1029c",
  1195 => x"d0ffc387",
  1196 => x"4bc0c84d",
  1197 => x"acb7c08c",
  1198 => x"c887c603",
  1199 => x"c04ba4c0",
  1200 => x"c4ccc44c",
  1201 => x"d049bf97",
  1202 => x"87d10299",
  1203 => x"ccc41ec0",
  1204 => x"ddff49cc",
  1205 => x"86c487db",
  1206 => x"ebc04a70",
  1207 => x"d0ffc387",
  1208 => x"ccccc41e",
  1209 => x"c8ddff49",
  1210 => x"7086c487",
  1211 => x"48d0ff4a",
  1212 => x"6e78c5c8",
  1213 => x"78d4c148",
  1214 => x"086e4815",
  1215 => x"058bc178",
  1216 => x"ff87f5ff",
  1217 => x"78c448d0",
  1218 => x"c5059a72",
  1219 => x"c148c087",
  1220 => x"1ec187cb",
  1221 => x"49ccccc4",
  1222 => x"87fadaff",
  1223 => x"9c7486c4",
  1224 => x"87c9fe05",
  1225 => x"c04866c4",
  1226 => x"d106a8b7",
  1227 => x"ccccc487",
  1228 => x"d078c048",
  1229 => x"f478c080",
  1230 => x"d8ccc480",
  1231 => x"66c478bf",
  1232 => x"a8b7c048",
  1233 => x"87d2fd01",
  1234 => x"d0ff4b6e",
  1235 => x"c178c548",
  1236 => x"7bc07bd3",
  1237 => x"48c178c4",
  1238 => x"c087c2c0",
  1239 => x"268ef448",
  1240 => x"264c264d",
  1241 => x"0e4f264b",
  1242 => x"5d5c5b5e",
  1243 => x"7186fc0e",
  1244 => x"4c4bc04d",
  1245 => x"e8c004ad",
  1246 => x"dec5c187",
  1247 => x"029c741e",
  1248 => x"4ac087c4",
  1249 => x"4ac187c2",
  1250 => x"e2e64972",
  1251 => x"7086c487",
  1252 => x"6e83c17e",
  1253 => x"7587c205",
  1254 => x"7584c14b",
  1255 => x"d8ff06ab",
  1256 => x"fc486e87",
  1257 => x"264d268e",
  1258 => x"264b264c",
  1259 => x"5b5e0e4f",
  1260 => x"fc0e5d5c",
  1261 => x"494c7186",
  1262 => x"cdc491de",
  1263 => x"85714de8",
  1264 => x"c1026d97",
  1265 => x"cdc487dd",
  1266 => x"7449bfd4",
  1267 => x"d6fe7181",
  1268 => x"487e7087",
  1269 => x"f3c00298",
  1270 => x"dccdc487",
  1271 => x"cb4a704b",
  1272 => x"ddf3fe49",
  1273 => x"cc4b7487",
  1274 => x"fcf3c193",
  1275 => x"c183c483",
  1276 => x"747bf0d0",
  1277 => x"dfc6c149",
  1278 => x"c17b7587",
  1279 => x"bf97e4f3",
  1280 => x"cdc41e49",
  1281 => x"d5c249dc",
  1282 => x"86c487ce",
  1283 => x"c6c14974",
  1284 => x"49c087c6",
  1285 => x"87e1c7c1",
  1286 => x"48c8ccc4",
  1287 => x"49c178c0",
  1288 => x"fc87c4de",
  1289 => x"264d268e",
  1290 => x"264b264c",
  1291 => x"0000004f",
  1292 => x"64616f4c",
  1293 => x"2e676e69",
  1294 => x"1e002e2e",
  1295 => x"4a711e73",
  1296 => x"d4cdc449",
  1297 => x"fc7181bf",
  1298 => x"4b7087dd",
  1299 => x"87c4029b",
  1300 => x"87e1e249",
  1301 => x"48d4cdc4",
  1302 => x"49c178c0",
  1303 => x"2687c8dd",
  1304 => x"1e4f264b",
  1305 => x"c6c149c0",
  1306 => x"4f2687cf",
  1307 => x"494a711e",
  1308 => x"f3c191cc",
  1309 => x"81c881fc",
  1310 => x"ccc44811",
  1311 => x"cdc458cc",
  1312 => x"78c048d4",
  1313 => x"dedc49c1",
  1314 => x"1e4f2687",
  1315 => x"d2029971",
  1316 => x"d8f5c187",
  1317 => x"f750c048",
  1318 => x"ecd1c180",
  1319 => x"f4f3c140",
  1320 => x"c187ce78",
  1321 => x"c148d4f5",
  1322 => x"fc78ecf3",
  1323 => x"e3d1c180",
  1324 => x"0e4f2678",
  1325 => x"5d5c5b5e",
  1326 => x"c386f40e",
  1327 => x"c04dd0ff",
  1328 => x"48a6c84c",
  1329 => x"7e7578c0",
  1330 => x"bfd4cdc4",
  1331 => x"06a8c048",
  1332 => x"c887c0c1",
  1333 => x"7e755ca6",
  1334 => x"48d0ffc3",
  1335 => x"f2c00298",
  1336 => x"4d66c487",
  1337 => x"1edec5c1",
  1338 => x"c40266cc",
  1339 => x"c24cc087",
  1340 => x"744cc187",
  1341 => x"87f7e049",
  1342 => x"7e7086c4",
  1343 => x"66c885c1",
  1344 => x"cc80c148",
  1345 => x"cdc458a6",
  1346 => x"03adbfd4",
  1347 => x"056e87c5",
  1348 => x"6e87d1ff",
  1349 => x"754cc04d",
  1350 => x"ddc3029d",
  1351 => x"dec5c187",
  1352 => x"0266cc1e",
  1353 => x"a6c887c7",
  1354 => x"c578c048",
  1355 => x"48a6c887",
  1356 => x"66c878c1",
  1357 => x"f6dfff49",
  1358 => x"7086c487",
  1359 => x"0298487e",
  1360 => x"4987e4c2",
  1361 => x"699781cb",
  1362 => x"0299d049",
  1363 => x"7487d4c1",
  1364 => x"c191cc49",
  1365 => x"c181fcf3",
  1366 => x"c879fbd0",
  1367 => x"51ffc381",
  1368 => x"91de4974",
  1369 => x"4de8cdc4",
  1370 => x"c1c28571",
  1371 => x"a5c17d97",
  1372 => x"51e0c049",
  1373 => x"97e0c7c4",
  1374 => x"87d202bf",
  1375 => x"a5c284c1",
  1376 => x"e0c7c44b",
  1377 => x"fe49db4a",
  1378 => x"c187f7ec",
  1379 => x"a5cd87d9",
  1380 => x"c151c049",
  1381 => x"4ba5c284",
  1382 => x"49cb4a6e",
  1383 => x"87e2ecfe",
  1384 => x"7487c4c1",
  1385 => x"c191cc49",
  1386 => x"c181fcf3",
  1387 => x"c479edce",
  1388 => x"bf97e0c7",
  1389 => x"7487d802",
  1390 => x"c191de49",
  1391 => x"e8cdc484",
  1392 => x"c483714b",
  1393 => x"dd4ae0c7",
  1394 => x"f5ebfe49",
  1395 => x"7487d887",
  1396 => x"c493de4b",
  1397 => x"cb83e8cd",
  1398 => x"51c049a3",
  1399 => x"6e7384c1",
  1400 => x"fe49cb4a",
  1401 => x"c887dbeb",
  1402 => x"80c14866",
  1403 => x"c758a6cc",
  1404 => x"c5c003ac",
  1405 => x"fc056e87",
  1406 => x"487487e3",
  1407 => x"4d268ef4",
  1408 => x"4b264c26",
  1409 => x"731e4f26",
  1410 => x"494b711e",
  1411 => x"f3c191cc",
  1412 => x"a1c881fc",
  1413 => x"e0f3c14a",
  1414 => x"c9501248",
  1415 => x"c8c14aa1",
  1416 => x"501248c4",
  1417 => x"f3c181ca",
  1418 => x"501148e4",
  1419 => x"97e4f3c1",
  1420 => x"c01e49bf",
  1421 => x"dfccc249",
  1422 => x"c8ccc487",
  1423 => x"c178de48",
  1424 => x"87e3d549",
  1425 => x"4b268efc",
  1426 => x"5e0e4f26",
  1427 => x"0e5d5c5b",
  1428 => x"4d7186f4",
  1429 => x"c191cc49",
  1430 => x"c881fcf3",
  1431 => x"a1ca4aa1",
  1432 => x"48a6c47e",
  1433 => x"bfe4d1c4",
  1434 => x"bf976e78",
  1435 => x"4c66c44b",
  1436 => x"48122c73",
  1437 => x"7058a6cc",
  1438 => x"c984c19c",
  1439 => x"49699781",
  1440 => x"c204acb7",
  1441 => x"6e4cc087",
  1442 => x"c84abf97",
  1443 => x"31724966",
  1444 => x"66c4b9ff",
  1445 => x"72487499",
  1446 => x"484a7030",
  1447 => x"d1c4b071",
  1448 => x"f9c158e8",
  1449 => x"49c087f1",
  1450 => x"7587fcd3",
  1451 => x"e7fbc049",
  1452 => x"268ef487",
  1453 => x"264c264d",
  1454 => x"1e4f264b",
  1455 => x"4b711e73",
  1456 => x"024aa3c6",
  1457 => x"8ac187db",
  1458 => x"8a87d602",
  1459 => x"87dac102",
  1460 => x"fcc0028a",
  1461 => x"c0028a87",
  1462 => x"028a87e1",
  1463 => x"dbc187cb",
  1464 => x"f649c787",
  1465 => x"dec187c6",
  1466 => x"d4cdc487",
  1467 => x"cbc102bf",
  1468 => x"88c14887",
  1469 => x"58d8cdc4",
  1470 => x"c487c1c1",
  1471 => x"02bfd8cd",
  1472 => x"c487f9c0",
  1473 => x"48bfd4cd",
  1474 => x"cdc480c1",
  1475 => x"ebc058d8",
  1476 => x"d4cdc487",
  1477 => x"89c649bf",
  1478 => x"59d8cdc4",
  1479 => x"03a9b7c0",
  1480 => x"cdc487da",
  1481 => x"78c048d4",
  1482 => x"cdc487d2",
  1483 => x"cb02bfd8",
  1484 => x"d4cdc487",
  1485 => x"80c648bf",
  1486 => x"58d8cdc4",
  1487 => x"e6d149c0",
  1488 => x"c0497387",
  1489 => x"2687d1f9",
  1490 => x"0e4f264b",
  1491 => x"5d5c5b5e",
  1492 => x"86d4ff0e",
  1493 => x"c859a6dc",
  1494 => x"78c048a6",
  1495 => x"c0c180c4",
  1496 => x"80c47866",
  1497 => x"80c478c1",
  1498 => x"cdc478c1",
  1499 => x"78c148d8",
  1500 => x"bfc8ccc4",
  1501 => x"05a8de48",
  1502 => x"f6f487c9",
  1503 => x"58a6cc87",
  1504 => x"c187dfcf",
  1505 => x"e487ecf7",
  1506 => x"f7c187e8",
  1507 => x"4c7087c2",
  1508 => x"02acfbc0",
  1509 => x"d887f0c1",
  1510 => x"e2c10566",
  1511 => x"66fcc087",
  1512 => x"6a82c44a",
  1513 => x"d8eec17e",
  1514 => x"20496e48",
  1515 => x"10412041",
  1516 => x"66fcc051",
  1517 => x"c6d8c148",
  1518 => x"c7496a78",
  1519 => x"c0517481",
  1520 => x"c84966fc",
  1521 => x"c051c181",
  1522 => x"c94966fc",
  1523 => x"c051c081",
  1524 => x"ca4966fc",
  1525 => x"c151c081",
  1526 => x"6a1ed81e",
  1527 => x"e381c849",
  1528 => x"86c887e5",
  1529 => x"4866c0c1",
  1530 => x"c701a8c0",
  1531 => x"48a6c887",
  1532 => x"87ce78c1",
  1533 => x"4866c0c1",
  1534 => x"a6d088c1",
  1535 => x"e287c358",
  1536 => x"a6d087f0",
  1537 => x"7478c248",
  1538 => x"d1cd029c",
  1539 => x"4866c887",
  1540 => x"a866c4c1",
  1541 => x"87c6cd03",
  1542 => x"c048a6dc",
  1543 => x"f4c17e78",
  1544 => x"4c7087ee",
  1545 => x"05acd0c1",
  1546 => x"c487d9c2",
  1547 => x"786e48a6",
  1548 => x"7087c1e4",
  1549 => x"d7f4c17e",
  1550 => x"c04c7087",
  1551 => x"c105acec",
  1552 => x"66c887ed",
  1553 => x"c091cc49",
  1554 => x"c48166fc",
  1555 => x"4d6a4aa1",
  1556 => x"6e4aa1c8",
  1557 => x"ecd1c152",
  1558 => x"f3f3c179",
  1559 => x"9c4c7087",
  1560 => x"c087d902",
  1561 => x"d302acfb",
  1562 => x"c1557487",
  1563 => x"7087e1f3",
  1564 => x"c7029c4c",
  1565 => x"acfbc087",
  1566 => x"87edff05",
  1567 => x"c255e0c0",
  1568 => x"97c055c1",
  1569 => x"4866d87d",
  1570 => x"05a866c4",
  1571 => x"66c887db",
  1572 => x"a866cc48",
  1573 => x"c887ca04",
  1574 => x"80c14866",
  1575 => x"c858a6cc",
  1576 => x"4866cc87",
  1577 => x"a6d088c1",
  1578 => x"e3f2c158",
  1579 => x"c14c7087",
  1580 => x"c805acd0",
  1581 => x"4866d487",
  1582 => x"a6d880c1",
  1583 => x"acd0c158",
  1584 => x"87e7fd02",
  1585 => x"66d8486e",
  1586 => x"e3c905a8",
  1587 => x"a6e0c087",
  1588 => x"7478c048",
  1589 => x"88fbc048",
  1590 => x"7058a6c8",
  1591 => x"e4c90298",
  1592 => x"88cb4887",
  1593 => x"7058a6c8",
  1594 => x"d1c10298",
  1595 => x"88c94887",
  1596 => x"7058a6c8",
  1597 => x"c1c40298",
  1598 => x"88c44887",
  1599 => x"7058a6c8",
  1600 => x"87cf0298",
  1601 => x"c888c148",
  1602 => x"987058a6",
  1603 => x"87eac302",
  1604 => x"dc87d4c8",
  1605 => x"f0c048a6",
  1606 => x"f3f0c178",
  1607 => x"c04c7087",
  1608 => x"c002acec",
  1609 => x"e0c087c4",
  1610 => x"ecc05ca6",
  1611 => x"cdc002ac",
  1612 => x"dbf0c187",
  1613 => x"c04c7087",
  1614 => x"ff05acec",
  1615 => x"ecc087f3",
  1616 => x"c4c002ac",
  1617 => x"c7f0c187",
  1618 => x"ca1ec087",
  1619 => x"4966d01e",
  1620 => x"c4c191cc",
  1621 => x"80714866",
  1622 => x"c858a6cc",
  1623 => x"80c44866",
  1624 => x"cc58a6d0",
  1625 => x"ff49bf66",
  1626 => x"c187dcdd",
  1627 => x"d41ede1e",
  1628 => x"ff49bf66",
  1629 => x"d087d0dd",
  1630 => x"48497086",
  1631 => x"c08808c0",
  1632 => x"c058a6e8",
  1633 => x"eec006a8",
  1634 => x"66e4c087",
  1635 => x"03a8dd48",
  1636 => x"c487e4c0",
  1637 => x"c049bf66",
  1638 => x"c08166e4",
  1639 => x"e4c051e0",
  1640 => x"81c14966",
  1641 => x"81bf66c4",
  1642 => x"c051c1c2",
  1643 => x"c24966e4",
  1644 => x"bf66c481",
  1645 => x"6e51c081",
  1646 => x"c6d8c148",
  1647 => x"c8496e78",
  1648 => x"5166d081",
  1649 => x"81c9496e",
  1650 => x"6e5166d4",
  1651 => x"dc81ca49",
  1652 => x"66d05166",
  1653 => x"d480c148",
  1654 => x"66c858a6",
  1655 => x"a866cc48",
  1656 => x"87cbc004",
  1657 => x"c14866c8",
  1658 => x"58a6cc80",
  1659 => x"cc87d6c5",
  1660 => x"88c14866",
  1661 => x"c558a6d0",
  1662 => x"dcff87cb",
  1663 => x"e8c087f6",
  1664 => x"dcff58a6",
  1665 => x"e0c087ee",
  1666 => x"ecc058a6",
  1667 => x"cac005a8",
  1668 => x"48a6dc87",
  1669 => x"7866e4c0",
  1670 => x"c187c4c0",
  1671 => x"c887f1ec",
  1672 => x"91cc4966",
  1673 => x"4866fcc0",
  1674 => x"a6c88071",
  1675 => x"4a66c458",
  1676 => x"66c482c8",
  1677 => x"c081ca49",
  1678 => x"dc5166e4",
  1679 => x"81c14966",
  1680 => x"8966e4c0",
  1681 => x"307148c1",
  1682 => x"89c14970",
  1683 => x"c47a9771",
  1684 => x"49bfe4d1",
  1685 => x"2966e4c0",
  1686 => x"484a6a97",
  1687 => x"ecc09871",
  1688 => x"66c458a6",
  1689 => x"6981c449",
  1690 => x"4866d84d",
  1691 => x"c002a86e",
  1692 => x"7ec087c5",
  1693 => x"c187c2c0",
  1694 => x"c01e6e7e",
  1695 => x"49751ee0",
  1696 => x"87c3d9ff",
  1697 => x"4c7086c8",
  1698 => x"06acb7c0",
  1699 => x"7487d0c1",
  1700 => x"49e0c085",
  1701 => x"4b758974",
  1702 => x"4ae4eec1",
  1703 => x"e1d8fe71",
  1704 => x"7585c287",
  1705 => x"66e0c07e",
  1706 => x"c080c148",
  1707 => x"c058a6e4",
  1708 => x"c14966e8",
  1709 => x"02a97081",
  1710 => x"c087c5c0",
  1711 => x"87c2c04d",
  1712 => x"1e754dc1",
  1713 => x"c049a4c2",
  1714 => x"887148e0",
  1715 => x"c81e4970",
  1716 => x"d7ff4966",
  1717 => x"86c887f1",
  1718 => x"01a8b7c0",
  1719 => x"c087c6ff",
  1720 => x"c00266e0",
  1721 => x"66c487d3",
  1722 => x"c081c949",
  1723 => x"c45166e0",
  1724 => x"d9c14866",
  1725 => x"cec078ca",
  1726 => x"4966c487",
  1727 => x"51c281c9",
  1728 => x"c34866c4",
  1729 => x"c878d0dd",
  1730 => x"66cc4866",
  1731 => x"cbc004a8",
  1732 => x"4866c887",
  1733 => x"a6cc80c1",
  1734 => x"87e9c058",
  1735 => x"c14866cc",
  1736 => x"58a6d088",
  1737 => x"ff87dec0",
  1738 => x"7087c7d6",
  1739 => x"87d5c04c",
  1740 => x"05acc6c1",
  1741 => x"d087c8c0",
  1742 => x"80c14866",
  1743 => x"ff58a6d4",
  1744 => x"7087efd5",
  1745 => x"4866d44c",
  1746 => x"a6d880c1",
  1747 => x"029c7458",
  1748 => x"c887cbc0",
  1749 => x"c4c14866",
  1750 => x"f204a866",
  1751 => x"d5ff87fa",
  1752 => x"66c887c7",
  1753 => x"03a8c748",
  1754 => x"c887e1c0",
  1755 => x"cdc44c66",
  1756 => x"78c048d8",
  1757 => x"91cc4974",
  1758 => x"8166fcc0",
  1759 => x"6a4aa1c4",
  1760 => x"7952c04a",
  1761 => x"acc784c1",
  1762 => x"87e2ff04",
  1763 => x"268ed4ff",
  1764 => x"264c264d",
  1765 => x"004f264b",
  1766 => x"64616f4c",
  1767 => x"202e2a20",
  1768 => x"00000000",
  1769 => x"1e00203a",
  1770 => x"4b711e73",
  1771 => x"87c6029b",
  1772 => x"48d4cdc4",
  1773 => x"1ec778c0",
  1774 => x"bfd4cdc4",
  1775 => x"fcf3c11e",
  1776 => x"c8ccc41e",
  1777 => x"c2ee49bf",
  1778 => x"c486cc87",
  1779 => x"49bfc8cc",
  1780 => x"7387f8e2",
  1781 => x"87c8029b",
  1782 => x"49fcf3c1",
  1783 => x"87c6e8c0",
  1784 => x"4f264b26",
  1785 => x"fc1e731e",
  1786 => x"4bffc386",
  1787 => x"fc4ad4ff",
  1788 => x"98c148bf",
  1789 => x"98487e70",
  1790 => x"87fbc002",
  1791 => x"c148d0ff",
  1792 => x"d2c278c1",
  1793 => x"c37a737a",
  1794 => x"4849d1ff",
  1795 => x"506a80ff",
  1796 => x"516a7a73",
  1797 => x"80c17a73",
  1798 => x"7a73506a",
  1799 => x"7a73506a",
  1800 => x"7a73496a",
  1801 => x"7a73506a",
  1802 => x"ffc3506a",
  1803 => x"ff5997da",
  1804 => x"c0c148d0",
  1805 => x"c387d778",
  1806 => x"4849d1ff",
  1807 => x"50c080ff",
  1808 => x"c080c151",
  1809 => x"c150d950",
  1810 => x"50e2c050",
  1811 => x"ffc350c3",
  1812 => x"50c048d7",
  1813 => x"8efc80f8",
  1814 => x"4f264b26",
  1815 => x"87d0cc1e",
  1816 => x"c2fd49c1",
  1817 => x"d1dcfe87",
  1818 => x"02987087",
  1819 => x"e5fe87cd",
  1820 => x"987087dd",
  1821 => x"c187c402",
  1822 => x"c087c24a",
  1823 => x"059a724a",
  1824 => x"1ec087ce",
  1825 => x"49f0f2c1",
  1826 => x"87e5f2c0",
  1827 => x"87fe86c4",
  1828 => x"f2c11ec0",
  1829 => x"f2c049fc",
  1830 => x"1ec087d7",
  1831 => x"87c2f9c1",
  1832 => x"f2c04970",
  1833 => x"d2c387cb",
  1834 => x"268ef887",
  1835 => x"0000004f",
  1836 => x"66204453",
  1837 => x"656c6961",
  1838 => x"00002e64",
  1839 => x"746f6f42",
  1840 => x"2e676e69",
  1841 => x"1e002e2e",
  1842 => x"48d4cdc4",
  1843 => x"ccc478c0",
  1844 => x"78c048c8",
  1845 => x"c187c5fe",
  1846 => x"c087e4fb",
  1847 => x"004f2648",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000001",
  1851 => x"78452080",
  1852 => x"00007469",
  1853 => x"61422080",
  1854 => x"00006b63",
  1855 => x"000013ad",
  1856 => x"00004368",
  1857 => x"00000000",
  1858 => x"000013ad",
  1859 => x"00004386",
  1860 => x"00000000",
  1861 => x"000013ad",
  1862 => x"000043a4",
  1863 => x"00000000",
  1864 => x"000013ad",
  1865 => x"000043c2",
  1866 => x"00000000",
  1867 => x"000013ad",
  1868 => x"000043e0",
  1869 => x"00000000",
  1870 => x"000013ad",
  1871 => x"000043fe",
  1872 => x"00000000",
  1873 => x"000013ad",
  1874 => x"0000441c",
  1875 => x"00000000",
  1876 => x"0000146c",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"000016bb",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"48f0fe1e",
  1883 => x"09cd78c0",
  1884 => x"4f260979",
  1885 => x"bff0fe1e",
  1886 => x"1e4f2648",
  1887 => x"c148f0fe",
  1888 => x"1e4f2678",
  1889 => x"c048f0fe",
  1890 => x"1e4f2678",
  1891 => x"97c04a71",
  1892 => x"49a2c17a",
  1893 => x"a2ca51c0",
  1894 => x"cb51c049",
  1895 => x"51c049a2",
  1896 => x"5e0e4f26",
  1897 => x"f00e5c5b",
  1898 => x"ca4c7186",
  1899 => x"699749a4",
  1900 => x"4ba4cb7e",
  1901 => x"c8486b97",
  1902 => x"80c158a6",
  1903 => x"c758a6cc",
  1904 => x"58a6d098",
  1905 => x"66cc486e",
  1906 => x"87db05a8",
  1907 => x"977e6997",
  1908 => x"a6c8486b",
  1909 => x"cc80c158",
  1910 => x"98c758a6",
  1911 => x"6e58a6d0",
  1912 => x"a866cc48",
  1913 => x"fe87e502",
  1914 => x"a4cc87d9",
  1915 => x"496b974a",
  1916 => x"dc49a172",
  1917 => x"6b975166",
  1918 => x"c1486e7e",
  1919 => x"58a6c880",
  1920 => x"a6cc98c7",
  1921 => x"7b977058",
  1922 => x"fd87d1c2",
  1923 => x"8ef087ed",
  1924 => x"4b264c26",
  1925 => x"5e0e4f26",
  1926 => x"0e5d5c5b",
  1927 => x"4d7186f4",
  1928 => x"c17e6d97",
  1929 => x"6c974ca5",
  1930 => x"58a6c848",
  1931 => x"66c4486e",
  1932 => x"87c505a8",
  1933 => x"e6c048ff",
  1934 => x"87c7fd87",
  1935 => x"9749a5c2",
  1936 => x"a3714b6c",
  1937 => x"4b6b974b",
  1938 => x"6e7e6c97",
  1939 => x"c880c148",
  1940 => x"98c758a6",
  1941 => x"7058a6cc",
  1942 => x"defc7c97",
  1943 => x"f4487387",
  1944 => x"264d268e",
  1945 => x"264b264c",
  1946 => x"5b5e0e4f",
  1947 => x"86f40e5c",
  1948 => x"66d84c71",
  1949 => x"9affc34a",
  1950 => x"974ba4c2",
  1951 => x"a173496c",
  1952 => x"97517249",
  1953 => x"486e7e6c",
  1954 => x"a6c880c1",
  1955 => x"cc98c758",
  1956 => x"547058a6",
  1957 => x"4c268ef4",
  1958 => x"4f264b26",
  1959 => x"f41e731e",
  1960 => x"87dffb86",
  1961 => x"494bbfe0",
  1962 => x"99c0e0c0",
  1963 => x"7387cb02",
  1964 => x"fcd0c41e",
  1965 => x"87f1fe49",
  1966 => x"497386c4",
  1967 => x"0299c0d0",
  1968 => x"c487c0c1",
  1969 => x"bf97c6d1",
  1970 => x"c7d1c47e",
  1971 => x"c848bf97",
  1972 => x"486e58a6",
  1973 => x"02a866c4",
  1974 => x"c487e8c0",
  1975 => x"bf97c6d1",
  1976 => x"c8d1c449",
  1977 => x"e0481181",
  1978 => x"d1c47808",
  1979 => x"7ebf97c6",
  1980 => x"80c1486e",
  1981 => x"c758a6c8",
  1982 => x"58a6cc98",
  1983 => x"48c6d1c4",
  1984 => x"e45066c8",
  1985 => x"c0494bbf",
  1986 => x"0299c0e0",
  1987 => x"1e7387cb",
  1988 => x"49d0d1c4",
  1989 => x"c487d2fd",
  1990 => x"d0497386",
  1991 => x"c10299c0",
  1992 => x"d1c487c0",
  1993 => x"7ebf97da",
  1994 => x"97dbd1c4",
  1995 => x"a6c848bf",
  1996 => x"c4486e58",
  1997 => x"c002a866",
  1998 => x"d1c487e8",
  1999 => x"49bf97da",
  2000 => x"81dcd1c4",
  2001 => x"08e44811",
  2002 => x"dad1c478",
  2003 => x"6e7ebf97",
  2004 => x"c880c148",
  2005 => x"98c758a6",
  2006 => x"c458a6cc",
  2007 => x"c848dad1",
  2008 => x"cff85066",
  2009 => x"f87e7087",
  2010 => x"8ef487d1",
  2011 => x"4f264b26",
  2012 => x"fcd0c41e",
  2013 => x"87d3f849",
  2014 => x"49d0d1c4",
  2015 => x"c187ccf8",
  2016 => x"f749dcfa",
  2017 => x"efc287e2",
  2018 => x"1e4f2687",
  2019 => x"d0c41e73",
  2020 => x"c1fa49fc",
  2021 => x"c04a7087",
  2022 => x"c204aab7",
  2023 => x"f0c387cc",
  2024 => x"87c905aa",
  2025 => x"48f0c0c2",
  2026 => x"edc178c1",
  2027 => x"aae0c387",
  2028 => x"c287c905",
  2029 => x"c148f4c0",
  2030 => x"87dec178",
  2031 => x"bff4c0c2",
  2032 => x"c287c602",
  2033 => x"c24ba2c0",
  2034 => x"c24b7287",
  2035 => x"02bff0c0",
  2036 => x"7387e0c0",
  2037 => x"29b7c449",
  2038 => x"ccc2c291",
  2039 => x"cf4a7381",
  2040 => x"c192c29a",
  2041 => x"70307248",
  2042 => x"72baff4a",
  2043 => x"70986948",
  2044 => x"7387db79",
  2045 => x"29b7c449",
  2046 => x"ccc2c291",
  2047 => x"cf4a7381",
  2048 => x"c392c29a",
  2049 => x"70307248",
  2050 => x"b069484a",
  2051 => x"c0c27970",
  2052 => x"78c048f4",
  2053 => x"48f0c0c2",
  2054 => x"d0c478c0",
  2055 => x"f5f749fc",
  2056 => x"c04a7087",
  2057 => x"fd03aab7",
  2058 => x"48c087f4",
  2059 => x"4f264b26",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"724ac01e",
  2063 => x"c291c449",
  2064 => x"c081ccc2",
  2065 => x"d082c179",
  2066 => x"ee04aab7",
  2067 => x"0e4f2687",
  2068 => x"5d5c5b5e",
  2069 => x"f44d710e",
  2070 => x"4a7587e9",
  2071 => x"922ab7c4",
  2072 => x"82ccc2c2",
  2073 => x"9ccf4c75",
  2074 => x"496a94c2",
  2075 => x"c32b744b",
  2076 => x"7448c29b",
  2077 => x"ff4c7030",
  2078 => x"714874bc",
  2079 => x"f37a7098",
  2080 => x"487387f9",
  2081 => x"4c264d26",
  2082 => x"4f264b26",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"48d0ff1e",
  2100 => x"7178e1c8",
  2101 => x"08d4ff48",
  2102 => x"1e4f2678",
  2103 => x"c848d0ff",
  2104 => x"487178e1",
  2105 => x"7808d4ff",
  2106 => x"ff4866c4",
  2107 => x"267808d4",
  2108 => x"4a711e4f",
  2109 => x"1e4966c4",
  2110 => x"deff4972",
  2111 => x"48d0ff87",
  2112 => x"fc78e0c0",
  2113 => x"1e4f268e",
  2114 => x"4b711e73",
  2115 => x"1e4966c8",
  2116 => x"e0c14a73",
  2117 => x"d8ff49a2",
  2118 => x"268efc87",
  2119 => x"1e4f264b",
  2120 => x"4b711e73",
  2121 => x"fe49e2c0",
  2122 => x"4ac787e2",
  2123 => x"d4ff4813",
  2124 => x"49727808",
  2125 => x"99718ac1",
  2126 => x"ff87f105",
  2127 => x"e0c048d0",
  2128 => x"264b2678",
  2129 => x"d0ff1e4f",
  2130 => x"78c9c848",
  2131 => x"d4ff4871",
  2132 => x"4f267808",
  2133 => x"494a711e",
  2134 => x"d0ff87eb",
  2135 => x"2678c848",
  2136 => x"1e731e4f",
  2137 => x"d1c44b71",
  2138 => x"c302bff4",
  2139 => x"87ebc287",
  2140 => x"c848d0ff",
  2141 => x"487378c9",
  2142 => x"ffb0e0c0",
  2143 => x"c47808d4",
  2144 => x"c048e8d1",
  2145 => x"0266c878",
  2146 => x"ffc387c5",
  2147 => x"c087c249",
  2148 => x"f0d1c449",
  2149 => x"0266cc59",
  2150 => x"d5c587c6",
  2151 => x"87c44ad5",
  2152 => x"4affffcf",
  2153 => x"5af4d1c4",
  2154 => x"48f4d1c4",
  2155 => x"4b2678c1",
  2156 => x"5e0e4f26",
  2157 => x"0e5d5c5b",
  2158 => x"d1c44d71",
  2159 => x"754bbff0",
  2160 => x"87cb029d",
  2161 => x"c291c849",
  2162 => x"714ad8c5",
  2163 => x"c287c482",
  2164 => x"c04ad8c9",
  2165 => x"7349124c",
  2166 => x"ecd1c499",
  2167 => x"b87148bf",
  2168 => x"7808d4ff",
  2169 => x"842bb7c1",
  2170 => x"04acb7c8",
  2171 => x"d1c487e7",
  2172 => x"c848bfe8",
  2173 => x"ecd1c480",
  2174 => x"264d2658",
  2175 => x"264b264c",
  2176 => x"1e731e4f",
  2177 => x"4a134b71",
  2178 => x"87cb029a",
  2179 => x"e1fe4972",
  2180 => x"9a4a1387",
  2181 => x"2687f505",
  2182 => x"1e4f264b",
  2183 => x"bfe8d1c4",
  2184 => x"e8d1c449",
  2185 => x"78a1c148",
  2186 => x"a9b7c0c4",
  2187 => x"ff87db03",
  2188 => x"d1c448d4",
  2189 => x"c478bfec",
  2190 => x"49bfe8d1",
  2191 => x"48e8d1c4",
  2192 => x"c478a1c1",
  2193 => x"04a9b7c0",
  2194 => x"d0ff87e5",
  2195 => x"c478c848",
  2196 => x"c048f4d1",
  2197 => x"004f2678",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"5f000000",
  2201 => x"0000005f",
  2202 => x"00030300",
  2203 => x"00000303",
  2204 => x"147f7f14",
  2205 => x"00147f7f",
  2206 => x"6b2e2400",
  2207 => x"00123a6b",
  2208 => x"18366a4c",
  2209 => x"0032566c",
  2210 => x"594f7e30",
  2211 => x"40683a77",
  2212 => x"07040000",
  2213 => x"00000003",
  2214 => x"3e1c0000",
  2215 => x"00004163",
  2216 => x"63410000",
  2217 => x"00001c3e",
  2218 => x"1c3e2a08",
  2219 => x"082a3e1c",
  2220 => x"3e080800",
  2221 => x"0008083e",
  2222 => x"e0800000",
  2223 => x"00000060",
  2224 => x"08080800",
  2225 => x"00080808",
  2226 => x"60000000",
  2227 => x"00000060",
  2228 => x"18306040",
  2229 => x"0103060c",
  2230 => x"597f3e00",
  2231 => x"003e7f4d",
  2232 => x"7f060400",
  2233 => x"0000007f",
  2234 => x"71634200",
  2235 => x"00464f59",
  2236 => x"49632200",
  2237 => x"00367f49",
  2238 => x"13161c18",
  2239 => x"00107f7f",
  2240 => x"45672700",
  2241 => x"00397d45",
  2242 => x"4b7e3c00",
  2243 => x"00307949",
  2244 => x"71010100",
  2245 => x"00070f79",
  2246 => x"497f3600",
  2247 => x"00367f49",
  2248 => x"494f0600",
  2249 => x"001e3f69",
  2250 => x"66000000",
  2251 => x"00000066",
  2252 => x"e6800000",
  2253 => x"00000066",
  2254 => x"14080800",
  2255 => x"00222214",
  2256 => x"14141400",
  2257 => x"00141414",
  2258 => x"14222200",
  2259 => x"00080814",
  2260 => x"51030200",
  2261 => x"00060f59",
  2262 => x"5d417f3e",
  2263 => x"001e1f55",
  2264 => x"097f7e00",
  2265 => x"007e7f09",
  2266 => x"497f7f00",
  2267 => x"00367f49",
  2268 => x"633e1c00",
  2269 => x"00414141",
  2270 => x"417f7f00",
  2271 => x"001c3e63",
  2272 => x"497f7f00",
  2273 => x"00414149",
  2274 => x"097f7f00",
  2275 => x"00010109",
  2276 => x"417f3e00",
  2277 => x"007a7b49",
  2278 => x"087f7f00",
  2279 => x"007f7f08",
  2280 => x"7f410000",
  2281 => x"0000417f",
  2282 => x"40602000",
  2283 => x"003f7f40",
  2284 => x"1c087f7f",
  2285 => x"00416336",
  2286 => x"407f7f00",
  2287 => x"00404040",
  2288 => x"0c067f7f",
  2289 => x"007f7f06",
  2290 => x"0c067f7f",
  2291 => x"007f7f18",
  2292 => x"417f3e00",
  2293 => x"003e7f41",
  2294 => x"097f7f00",
  2295 => x"00060f09",
  2296 => x"61417f3e",
  2297 => x"00407e7f",
  2298 => x"097f7f00",
  2299 => x"00667f19",
  2300 => x"4d6f2600",
  2301 => x"00327b59",
  2302 => x"7f010100",
  2303 => x"0001017f",
  2304 => x"407f3f00",
  2305 => x"003f7f40",
  2306 => x"703f0f00",
  2307 => x"000f3f70",
  2308 => x"18307f7f",
  2309 => x"007f7f30",
  2310 => x"1c366341",
  2311 => x"4163361c",
  2312 => x"7c060301",
  2313 => x"0103067c",
  2314 => x"4d597161",
  2315 => x"00414347",
  2316 => x"7f7f0000",
  2317 => x"00004141",
  2318 => x"0c060301",
  2319 => x"40603018",
  2320 => x"41410000",
  2321 => x"00007f7f",
  2322 => x"03060c08",
  2323 => x"00080c06",
  2324 => x"80808080",
  2325 => x"00808080",
  2326 => x"03000000",
  2327 => x"00000407",
  2328 => x"54742000",
  2329 => x"00787c54",
  2330 => x"447f7f00",
  2331 => x"00387c44",
  2332 => x"447c3800",
  2333 => x"00004444",
  2334 => x"447c3800",
  2335 => x"007f7f44",
  2336 => x"547c3800",
  2337 => x"00185c54",
  2338 => x"7f7e0400",
  2339 => x"00000505",
  2340 => x"a4bc1800",
  2341 => x"007cfca4",
  2342 => x"047f7f00",
  2343 => x"00787c04",
  2344 => x"3d000000",
  2345 => x"0000407d",
  2346 => x"80808000",
  2347 => x"00007dfd",
  2348 => x"107f7f00",
  2349 => x"00446c38",
  2350 => x"3f000000",
  2351 => x"0000407f",
  2352 => x"180c7c7c",
  2353 => x"00787c0c",
  2354 => x"047c7c00",
  2355 => x"00787c04",
  2356 => x"447c3800",
  2357 => x"00387c44",
  2358 => x"24fcfc00",
  2359 => x"00183c24",
  2360 => x"243c1800",
  2361 => x"00fcfc24",
  2362 => x"047c7c00",
  2363 => x"00080c04",
  2364 => x"545c4800",
  2365 => x"00207454",
  2366 => x"7f3f0400",
  2367 => x"00004444",
  2368 => x"407c3c00",
  2369 => x"007c7c40",
  2370 => x"603c1c00",
  2371 => x"001c3c60",
  2372 => x"30607c3c",
  2373 => x"003c7c60",
  2374 => x"10386c44",
  2375 => x"00446c38",
  2376 => x"e0bc1c00",
  2377 => x"001c3c60",
  2378 => x"74644400",
  2379 => x"00444c5c",
  2380 => x"3e080800",
  2381 => x"00414177",
  2382 => x"7f000000",
  2383 => x"0000007f",
  2384 => x"77414100",
  2385 => x"0008083e",
  2386 => x"03010102",
  2387 => x"00010202",
  2388 => x"7f7f7f7f",
  2389 => x"007f7f7f",
  2390 => x"1c1c0808",
  2391 => x"7f7f3e3e",
  2392 => x"3e3e7f7f",
  2393 => x"08081c1c",
  2394 => x"7c181000",
  2395 => x"0010187c",
  2396 => x"7c301000",
  2397 => x"0010307c",
  2398 => x"60603010",
  2399 => x"00061e78",
  2400 => x"183c6642",
  2401 => x"0042663c",
  2402 => x"c26a3878",
  2403 => x"00386cc6",
  2404 => x"60000060",
  2405 => x"00600000",
  2406 => x"5c5b5e0e",
  2407 => x"86fc0e5d",
  2408 => x"d2c47e71",
  2409 => x"c04cbfc8",
  2410 => x"c41ec04b",
  2411 => x"c402ab66",
  2412 => x"c24dc087",
  2413 => x"754dc187",
  2414 => x"ee49731e",
  2415 => x"86c887e3",
  2416 => x"ef49e0c0",
  2417 => x"a4c487ec",
  2418 => x"f0496a4a",
  2419 => x"caf187f3",
  2420 => x"c184cc87",
  2421 => x"abb7c883",
  2422 => x"87cdff04",
  2423 => x"4d268efc",
  2424 => x"4b264c26",
  2425 => x"711e4f26",
  2426 => x"ccd2c44a",
  2427 => x"ccd2c45a",
  2428 => x"4978c748",
  2429 => x"2687e1fe",
  2430 => x"1e731e4f",
  2431 => x"b7c04a71",
  2432 => x"87d303aa",
  2433 => x"bfd4e6c2",
  2434 => x"c187c405",
  2435 => x"c087c24b",
  2436 => x"d8e6c24b",
  2437 => x"c287c45b",
  2438 => x"c25ad8e6",
  2439 => x"4abfd4e6",
  2440 => x"c0c19ac1",
  2441 => x"ebec49a2",
  2442 => x"c248fc87",
  2443 => x"78bfd4e6",
  2444 => x"4f264b26",
  2445 => x"d4e6c21e",
  2446 => x"4f2648bf",
  2447 => x"c44a711e",
  2448 => x"49721e66",
  2449 => x"fc87c0eb",
  2450 => x"1e4f268e",
  2451 => x"c348d4ff",
  2452 => x"d0ff78ff",
  2453 => x"78e1c048",
  2454 => x"c148d4ff",
  2455 => x"c4487178",
  2456 => x"08d4ff30",
  2457 => x"48d0ff78",
  2458 => x"2678e0c0",
  2459 => x"e6c21e4f",
  2460 => x"c149bfd4",
  2461 => x"c487f5d4",
  2462 => x"e848c0d2",
  2463 => x"d1c478bf",
  2464 => x"bfec48fc",
  2465 => x"c0d2c478",
  2466 => x"c3494abf",
  2467 => x"b7c899ff",
  2468 => x"7148722a",
  2469 => x"c8d2c4b0",
  2470 => x"0e4f2658",
  2471 => x"5d5c5b5e",
  2472 => x"ff4b710e",
  2473 => x"d1c487c7",
  2474 => x"50c048f8",
  2475 => x"dee64973",
  2476 => x"4c497087",
  2477 => x"eecb9cc2",
  2478 => x"87e0cb49",
  2479 => x"d1c44d70",
  2480 => x"05bf97f8",
  2481 => x"d087e2c1",
  2482 => x"d2c44966",
  2483 => x"0599bfc4",
  2484 => x"66d487d6",
  2485 => x"fcd1c449",
  2486 => x"cb0599bf",
  2487 => x"e5497387",
  2488 => x"987087ed",
  2489 => x"87c1c102",
  2490 => x"c0fe4cc1",
  2491 => x"ca497587",
  2492 => x"987087f6",
  2493 => x"c487c602",
  2494 => x"c148f8d1",
  2495 => x"f8d1c450",
  2496 => x"c005bf97",
  2497 => x"d2c487e3",
  2498 => x"d049bfc4",
  2499 => x"ff059966",
  2500 => x"d1c487d6",
  2501 => x"d449bffc",
  2502 => x"ff059966",
  2503 => x"497387ca",
  2504 => x"7087ece4",
  2505 => x"fffe0598",
  2506 => x"26487487",
  2507 => x"264c264d",
  2508 => x"0e4f264b",
  2509 => x"5d5c5b5e",
  2510 => x"c086f80e",
  2511 => x"bfec4c4d",
  2512 => x"48a6c47e",
  2513 => x"bfc8d2c4",
  2514 => x"c01ec178",
  2515 => x"fd49c71e",
  2516 => x"86c887c9",
  2517 => x"cd029870",
  2518 => x"fa49ff87",
  2519 => x"dac187db",
  2520 => x"87ebe349",
  2521 => x"d1c44dc1",
  2522 => x"02bf97f8",
  2523 => x"e6c287cf",
  2524 => x"c149bfcc",
  2525 => x"d0e6c2b9",
  2526 => x"cefb7159",
  2527 => x"c0d2c487",
  2528 => x"e6c24bbf",
  2529 => x"c005bfd4",
  2530 => x"fdc387e9",
  2531 => x"87ffe249",
  2532 => x"e249fac3",
  2533 => x"497387f9",
  2534 => x"7199ffc3",
  2535 => x"fa49c01e",
  2536 => x"497387da",
  2537 => x"7129b7c8",
  2538 => x"fa49c11e",
  2539 => x"86c887ce",
  2540 => x"c487f4c5",
  2541 => x"4bbfc4d2",
  2542 => x"87dd029b",
  2543 => x"bfd0e6c2",
  2544 => x"87e4c749",
  2545 => x"c4059870",
  2546 => x"d24bc087",
  2547 => x"49e0c287",
  2548 => x"c287c9c7",
  2549 => x"c658d4e6",
  2550 => x"d0e6c287",
  2551 => x"7378c048",
  2552 => x"0599c249",
  2553 => x"ebc387cd",
  2554 => x"87e3e149",
  2555 => x"99c24970",
  2556 => x"fb87c202",
  2557 => x"c149734c",
  2558 => x"87cd0599",
  2559 => x"e149f4c3",
  2560 => x"497087cd",
  2561 => x"c20299c2",
  2562 => x"734cfa87",
  2563 => x"0599c849",
  2564 => x"f5c387cd",
  2565 => x"87f7e049",
  2566 => x"99c24970",
  2567 => x"c487d502",
  2568 => x"02bfccd2",
  2569 => x"c14887ca",
  2570 => x"d0d2c488",
  2571 => x"87c2c058",
  2572 => x"4dc14cff",
  2573 => x"99c44973",
  2574 => x"c387cd05",
  2575 => x"cee049f2",
  2576 => x"c2497087",
  2577 => x"87dc0299",
  2578 => x"bfccd2c4",
  2579 => x"b7c7487e",
  2580 => x"cbc003a8",
  2581 => x"c1486e87",
  2582 => x"d0d2c480",
  2583 => x"87c2c058",
  2584 => x"4dc14cfe",
  2585 => x"ff49fdc3",
  2586 => x"7087e4df",
  2587 => x"0299c249",
  2588 => x"d2c487d5",
  2589 => x"c002bfcc",
  2590 => x"d2c487c9",
  2591 => x"78c048cc",
  2592 => x"fd87c2c0",
  2593 => x"c34dc14c",
  2594 => x"dfff49fa",
  2595 => x"497087c1",
  2596 => x"c00299c2",
  2597 => x"d2c487d9",
  2598 => x"c748bfcc",
  2599 => x"c003a8b7",
  2600 => x"d2c487c9",
  2601 => x"78c748cc",
  2602 => x"fc87c2c0",
  2603 => x"c04dc14c",
  2604 => x"c003acb7",
  2605 => x"66c487d3",
  2606 => x"80e0c148",
  2607 => x"bf6e7e70",
  2608 => x"87c5c002",
  2609 => x"7349744b",
  2610 => x"c31ec00f",
  2611 => x"dac11ef0",
  2612 => x"87c7f749",
  2613 => x"987086c8",
  2614 => x"87d8c002",
  2615 => x"bfccd2c4",
  2616 => x"cc496e7e",
  2617 => x"4a66c491",
  2618 => x"026a8271",
  2619 => x"4b87c5c0",
  2620 => x"0f73496e",
  2621 => x"c0029d75",
  2622 => x"d2c487c8",
  2623 => x"f249bfcc",
  2624 => x"e6c287d6",
  2625 => x"c002bfd8",
  2626 => x"c24987dd",
  2627 => x"987087da",
  2628 => x"87d3c002",
  2629 => x"bfccd2c4",
  2630 => x"87fcf149",
  2631 => x"d8f349c0",
  2632 => x"d8e6c287",
  2633 => x"f878c048",
  2634 => x"264d268e",
  2635 => x"264b264c",
  2636 => x"5b5e0e4f",
  2637 => x"fc0e5d5c",
  2638 => x"c44c7186",
  2639 => x"49bfc8d2",
  2640 => x"4da1d4c1",
  2641 => x"6981d8c1",
  2642 => x"029c747e",
  2643 => x"a5c487cf",
  2644 => x"c47b744b",
  2645 => x"49bfc8d2",
  2646 => x"6e87cbf2",
  2647 => x"059c747b",
  2648 => x"4bc087c4",
  2649 => x"4bc187c2",
  2650 => x"ccf24973",
  2651 => x"0266d487",
  2652 => x"c04987c8",
  2653 => x"4a7087e6",
  2654 => x"4ac087c2",
  2655 => x"5adce6c2",
  2656 => x"4d268efc",
  2657 => x"4b264c26",
  2658 => x"00004f26",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"ff4a711e",
  2664 => x"7249bfc8",
  2665 => x"4f2648a1",
  2666 => x"bfc8ff1e",
  2667 => x"c0c0fe89",
  2668 => x"a9c0c0c0",
  2669 => x"c087c401",
  2670 => x"c187c24a",
  2671 => x"2648724a",
  2672 => x"5b5e0e4f",
  2673 => x"710e5d5c",
  2674 => x"4cd4ff4b",
  2675 => x"c04866d0",
  2676 => x"ff49d678",
  2677 => x"c387f5db",
  2678 => x"496c7cff",
  2679 => x"7199ffc3",
  2680 => x"f0c3494d",
  2681 => x"a9e0c199",
  2682 => x"c387cb05",
  2683 => x"486c7cff",
  2684 => x"66d098c3",
  2685 => x"ffc37808",
  2686 => x"494a6c7c",
  2687 => x"ffc331c8",
  2688 => x"714a6c7c",
  2689 => x"c84972b2",
  2690 => x"7cffc331",
  2691 => x"b2714a6c",
  2692 => x"31c84972",
  2693 => x"6c7cffc3",
  2694 => x"ffb2714a",
  2695 => x"e0c048d0",
  2696 => x"029b7378",
  2697 => x"7b7287c2",
  2698 => x"4d264875",
  2699 => x"4b264c26",
  2700 => x"261e4f26",
  2701 => x"5b5e0e4f",
  2702 => x"86f80e5c",
  2703 => x"a6c81e76",
  2704 => x"87fdfd49",
  2705 => x"4b7086c4",
  2706 => x"a8c4486e",
  2707 => x"87f4c203",
  2708 => x"f0c34a73",
  2709 => x"aad0c19a",
  2710 => x"c187c702",
  2711 => x"c205aae0",
  2712 => x"497387e2",
  2713 => x"c30299c8",
  2714 => x"87c6ff87",
  2715 => x"9cc34c73",
  2716 => x"c105acc2",
  2717 => x"66c487c4",
  2718 => x"7131c949",
  2719 => x"4a66c41e",
  2720 => x"c492c8c1",
  2721 => x"7249d0d2",
  2722 => x"fec3fe81",
  2723 => x"ff49d887",
  2724 => x"c887f9d8",
  2725 => x"ffc31ec0",
  2726 => x"dbfd49d0",
  2727 => x"d0ff87c9",
  2728 => x"78e0c048",
  2729 => x"1ed0ffc3",
  2730 => x"c14a66cc",
  2731 => x"d2c492c8",
  2732 => x"817249d0",
  2733 => x"87c8fffd",
  2734 => x"acc186cc",
  2735 => x"87c4c105",
  2736 => x"c94966c4",
  2737 => x"c41e7131",
  2738 => x"c8c14a66",
  2739 => x"d0d2c492",
  2740 => x"fe817249",
  2741 => x"c387f4c2",
  2742 => x"c81ed0ff",
  2743 => x"c8c14a66",
  2744 => x"d0d2c492",
  2745 => x"fd817249",
  2746 => x"d787c6fd",
  2747 => x"dbd7ff49",
  2748 => x"1ec0c887",
  2749 => x"49d0ffc3",
  2750 => x"87c8d9fd",
  2751 => x"d0ff86cc",
  2752 => x"78e0c048",
  2753 => x"4c268ef8",
  2754 => x"4f264b26",
  2755 => x"5c5b5e0e",
  2756 => x"4a710e5d",
  2757 => x"d04cd4ff",
  2758 => x"b7c34d66",
  2759 => x"87c506ad",
  2760 => x"e2c148c0",
  2761 => x"751e7287",
  2762 => x"93c8c14b",
  2763 => x"83d0d2c4",
  2764 => x"f5fd4973",
  2765 => x"83c887fd",
  2766 => x"d0ff4b6b",
  2767 => x"78e1c848",
  2768 => x"48737cdd",
  2769 => x"7098ffc3",
  2770 => x"c849737c",
  2771 => x"487129b7",
  2772 => x"7098ffc3",
  2773 => x"d049737c",
  2774 => x"487129b7",
  2775 => x"7098ffc3",
  2776 => x"d848737c",
  2777 => x"7c7028b7",
  2778 => x"7c7c7cc0",
  2779 => x"7c7c7c7c",
  2780 => x"7c7c7c7c",
  2781 => x"48d0ff7c",
  2782 => x"7578e0c0",
  2783 => x"ff49dc1e",
  2784 => x"c887eed5",
  2785 => x"26487386",
  2786 => x"264c264d",
  2787 => x"1e4f264b",
  2788 => x"86fc1e73",
  2789 => x"f0c04b71",
  2790 => x"ecc04aa3",
  2791 => x"826949a3",
  2792 => x"695266cc",
  2793 => x"7080c148",
  2794 => x"98cf487e",
  2795 => x"8efc7970",
  2796 => x"4f264b26",
  2797 => x"5c5b5e0e",
  2798 => x"e94b710e",
  2799 => x"4c7087f6",
  2800 => x"87ffc6ff",
  2801 => x"c24966cc",
  2802 => x"dc0299c0",
  2803 => x"059c7487",
  2804 => x"e0c387ca",
  2805 => x"fe49731e",
  2806 => x"86c487f5",
  2807 => x"c41ee0c3",
  2808 => x"ff49fcd0",
  2809 => x"c487c2ca",
  2810 => x"4966cc86",
  2811 => x"0299c0c4",
  2812 => x"9c7487dc",
  2813 => x"c387ca05",
  2814 => x"49731ef0",
  2815 => x"c487d0fe",
  2816 => x"1ef0c386",
  2817 => x"49fcd0c4",
  2818 => x"87ddc9ff",
  2819 => x"9c7486c4",
  2820 => x"cc87cf05",
  2821 => x"ffc14966",
  2822 => x"731e7199",
  2823 => x"87effd49",
  2824 => x"66cc86c4",
  2825 => x"99ffc149",
  2826 => x"d0c41e71",
  2827 => x"c8ff49fc",
  2828 => x"c5ff87f7",
  2829 => x"8efc87c5",
  2830 => x"4b264c26",
  2831 => x"5e0e4f26",
  2832 => x"fc0e5c5b",
  2833 => x"fac4ff86",
  2834 => x"c0f3c287",
  2835 => x"d7f549bf",
  2836 => x"02987087",
  2837 => x"c487dcc1",
  2838 => x"48bfdcd7",
  2839 => x"bfe0d7c4",
  2840 => x"cec102a8",
  2841 => x"e4d7c487",
  2842 => x"dcd7c449",
  2843 => x"4c1181bf",
  2844 => x"aae0c34a",
  2845 => x"c387c602",
  2846 => x"c405aaf0",
  2847 => x"c24bc487",
  2848 => x"734bcf87",
  2849 => x"87d4f449",
  2850 => x"58c4f3c2",
  2851 => x"c848d0ff",
  2852 => x"d4ff78e1",
  2853 => x"7478c548",
  2854 => x"08d4ff48",
  2855 => x"48d0ff78",
  2856 => x"c478e0c0",
  2857 => x"48bfdcd7",
  2858 => x"7e7080c1",
  2859 => x"c498cf48",
  2860 => x"ff58e0d7",
  2861 => x"fc87c4c3",
  2862 => x"264c268e",
  2863 => x"004f264b",
  2864 => x"00000000",
  2865 => x"5c5b5e0e",
  2866 => x"dcff0e5d",
  2867 => x"c47ec086",
  2868 => x"49bff8d6",
  2869 => x"1e7181c2",
  2870 => x"4ac61e72",
  2871 => x"87f3d0fd",
  2872 => x"4a264871",
  2873 => x"a6cc4926",
  2874 => x"f8d6c458",
  2875 => x"81c449bf",
  2876 => x"1e721e71",
  2877 => x"d0fd4ac6",
  2878 => x"487187d9",
  2879 => x"49264a26",
  2880 => x"fc58a6d0",
  2881 => x"fec287f8",
  2882 => x"f249bfd4",
  2883 => x"987087da",
  2884 => x"87f4c902",
  2885 => x"f249e0c0",
  2886 => x"fec287c2",
  2887 => x"4cc058d8",
  2888 => x"91c44974",
  2889 => x"6981d0fe",
  2890 => x"c449744a",
  2891 => x"81bff8d6",
  2892 => x"d7c491c4",
  2893 => x"797281c4",
  2894 => x"87d2029a",
  2895 => x"89c14972",
  2896 => x"486e9a71",
  2897 => x"7e7080c1",
  2898 => x"ff059a72",
  2899 => x"84c187ee",
  2900 => x"04acb7c2",
  2901 => x"6e87c9ff",
  2902 => x"b7fcc048",
  2903 => x"e7c804a8",
  2904 => x"744cc087",
  2905 => x"8266c84a",
  2906 => x"d7c492c4",
  2907 => x"497482c4",
  2908 => x"c48166cc",
  2909 => x"c4d7c491",
  2910 => x"694a6a81",
  2911 => x"74b97249",
  2912 => x"f8d6c44b",
  2913 => x"93c483bf",
  2914 => x"83c4d7c4",
  2915 => x"4872ba6b",
  2916 => x"a6d89871",
  2917 => x"c4497458",
  2918 => x"81bff8d6",
  2919 => x"d7c491c4",
  2920 => x"7e6981c4",
  2921 => x"c048a6d8",
  2922 => x"5ca6d478",
  2923 => x"df4966d4",
  2924 => x"e2c60229",
  2925 => x"4a66d087",
  2926 => x"d892e0c0",
  2927 => x"ffc08266",
  2928 => x"70887248",
  2929 => x"48a6dc4a",
  2930 => x"80c478c0",
  2931 => x"496e78c0",
  2932 => x"4c7129df",
  2933 => x"48f4d6c4",
  2934 => x"497278c1",
  2935 => x"2ab731c3",
  2936 => x"ffc0b172",
  2937 => x"c391c499",
  2938 => x"714dc8f0",
  2939 => x"494b6d85",
  2940 => x"99c0c0c4",
  2941 => x"7487d602",
  2942 => x"c7c0029c",
  2943 => x"c080c887",
  2944 => x"87d3c578",
  2945 => x"48fcd6c4",
  2946 => x"cac578c1",
  2947 => x"029c7487",
  2948 => x"497387d8",
  2949 => x"99c0c0c2",
  2950 => x"87c3c002",
  2951 => x"6d2bb7d0",
  2952 => x"fffffd48",
  2953 => x"c07d7098",
  2954 => x"d6c487f8",
  2955 => x"c002bffc",
  2956 => x"487387f0",
  2957 => x"c828b7d0",
  2958 => x"987058a6",
  2959 => x"87e2c002",
  2960 => x"bfc0d7c4",
  2961 => x"c0e0c049",
  2962 => x"cac00299",
  2963 => x"c0497087",
  2964 => x"0299c0e0",
  2965 => x"6d87cbc0",
  2966 => x"c0c0c248",
  2967 => x"c47d70b0",
  2968 => x"49734b66",
  2969 => x"99c0c0c8",
  2970 => x"87c9c202",
  2971 => x"bfc0d7c4",
  2972 => x"9ac0cc4a",
  2973 => x"87cfc002",
  2974 => x"028ac0c4",
  2975 => x"8a87d8c0",
  2976 => x"87fac002",
  2977 => x"7387dfc1",
  2978 => x"99ffc349",
  2979 => x"efc391c2",
  2980 => x"4b1181fc",
  2981 => x"7387dec1",
  2982 => x"99ffc349",
  2983 => x"efc391c2",
  2984 => x"81c181fc",
  2985 => x"9c744b11",
  2986 => x"87c9c002",
  2987 => x"48a6e0c0",
  2988 => x"c0c178d2",
  2989 => x"48a6dc87",
  2990 => x"c078d2c4",
  2991 => x"497387f7",
  2992 => x"c299ffc3",
  2993 => x"fcefc391",
  2994 => x"1181c181",
  2995 => x"029c744b",
  2996 => x"c087cac0",
  2997 => x"c148a6e0",
  2998 => x"d8c078d9",
  2999 => x"48a6dc87",
  3000 => x"c078d9c5",
  3001 => x"497387cf",
  3002 => x"c299ffc3",
  3003 => x"fcefc391",
  3004 => x"1181c181",
  3005 => x"029c744b",
  3006 => x"7387dcc0",
  3007 => x"c7b9ff49",
  3008 => x"7199c0fc",
  3009 => x"c0d7c448",
  3010 => x"d7c498bf",
  3011 => x"ffc358c4",
  3012 => x"b3c0c49b",
  3013 => x"7387d4c0",
  3014 => x"c0fcc749",
  3015 => x"c4487199",
  3016 => x"b0bfc0d7",
  3017 => x"58c4d7c4",
  3018 => x"dc9bffc3",
  3019 => x"cac00266",
  3020 => x"d6c41e87",
  3021 => x"fbf149f4",
  3022 => x"7386c487",
  3023 => x"f4d6c41e",
  3024 => x"87f0f149",
  3025 => x"e0c086c4",
  3026 => x"cac00266",
  3027 => x"d6c41e87",
  3028 => x"dff149f4",
  3029 => x"d486c487",
  3030 => x"30c14866",
  3031 => x"6e58a6d8",
  3032 => x"7030c148",
  3033 => x"4866d87e",
  3034 => x"a6dc80c1",
  3035 => x"b7e0c058",
  3036 => x"f7f804a8",
  3037 => x"4c66d087",
  3038 => x"b7c284c1",
  3039 => x"e2f704ac",
  3040 => x"f8d6c487",
  3041 => x"7866c848",
  3042 => x"268edcff",
  3043 => x"264c264d",
  3044 => x"004f264b",
  3045 => x"00000000",
  3046 => x"724ac01e",
  3047 => x"c491c449",
  3048 => x"ff81c4d7",
  3049 => x"c682c179",
  3050 => x"ee04aab7",
  3051 => x"f8d6c487",
  3052 => x"4040c048",
  3053 => x"0e4f2678",
  3054 => x"0e5c5b5e",
  3055 => x"d4ff4a71",
  3056 => x"4b66cc4c",
  3057 => x"c848d0ff",
  3058 => x"7cc278c5",
  3059 => x"8bc14973",
  3060 => x"cd029971",
  3061 => x"127c1287",
  3062 => x"c149737c",
  3063 => x"0599718b",
  3064 => x"d0ff87f3",
  3065 => x"2678c448",
  3066 => x"264b264c",
  3067 => x"4a711e4f",
  3068 => x"c848d0ff",
  3069 => x"d4ff78c5",
  3070 => x"c878c348",
  3071 => x"49721ec0",
  3072 => x"87e3c5fd",
  3073 => x"c448d0ff",
  3074 => x"268efc78",
  3075 => x"d0ff1e4f",
  3076 => x"78c5c848",
  3077 => x"c648d4ff",
  3078 => x"ff487178",
  3079 => x"ff7808d4",
  3080 => x"78c448d0",
  3081 => x"ff1e4f26",
  3082 => x"c5c848d0",
  3083 => x"48d4ff78",
  3084 => x"d0ff78ca",
  3085 => x"2678c448",
  3086 => x"5b5e0e4f",
  3087 => x"ff0e5d5c",
  3088 => x"7e7186d4",
  3089 => x"81ca496e",
  3090 => x"48496997",
  3091 => x"d428b7c5",
  3092 => x"496e58a6",
  3093 => x"699781c1",
  3094 => x"b7c54849",
  3095 => x"58a6d828",
  3096 => x"48bf976e",
  3097 => x"df58a6dc",
  3098 => x"c0c0d099",
  3099 => x"c24a6e91",
  3100 => x"c0481282",
  3101 => x"7058a6e0",
  3102 => x"92c0c44a",
  3103 => x"6e49a172",
  3104 => x"1282c34a",
  3105 => x"a6e4c048",
  3106 => x"c0817058",
  3107 => x"6e59a6e8",
  3108 => x"c880c448",
  3109 => x"66c458a6",
  3110 => x"9c4cbf97",
  3111 => x"c487c305",
  3112 => x"66d04cc0",
  3113 => x"a8b7c248",
  3114 => x"87f1cf03",
  3115 => x"c14966d0",
  3116 => x"d4c491c8",
  3117 => x"807148e0",
  3118 => x"cc58a6d0",
  3119 => x"80c84866",
  3120 => x"c858a6cc",
  3121 => x"cf02bf66",
  3122 => x"c94887d3",
  3123 => x"a6ecc028",
  3124 => x"0266d858",
  3125 => x"4d87e3c2",
  3126 => x"c3028dc3",
  3127 => x"8dc187c3",
  3128 => x"87d6c202",
  3129 => x"c4028dc4",
  3130 => x"8dc287cf",
  3131 => x"87d6c702",
  3132 => x"ca028dc8",
  3133 => x"028d87e5",
  3134 => x"cb87e6cc",
  3135 => x"87cf028d",
  3136 => x"c3028dc3",
  3137 => x"8dc287f3",
  3138 => x"87fac602",
  3139 => x"d487fccd",
  3140 => x"d3c10566",
  3141 => x"d0ffc387",
  3142 => x"c84ac04b",
  3143 => x"fefc49c0",
  3144 => x"e8c087f0",
  3145 => x"89c14966",
  3146 => x"2ad84a71",
  3147 => x"97d4ffc3",
  3148 => x"d04a715a",
  3149 => x"d5ffc32a",
  3150 => x"4a715a97",
  3151 => x"ffc32ac8",
  3152 => x"c35a97d6",
  3153 => x"5997d7ff",
  3154 => x"c280c348",
  3155 => x"f91ec450",
  3156 => x"e2f949a0",
  3157 => x"c086c487",
  3158 => x"87f1fa49",
  3159 => x"49e0d3c3",
  3160 => x"c08166d0",
  3161 => x"87f8cc51",
  3162 => x"e0fa49c2",
  3163 => x"e0d3c387",
  3164 => x"8166d049",
  3165 => x"cc51e5c0",
  3166 => x"66d487e6",
  3167 => x"c387d005",
  3168 => x"d049e0d3",
  3169 => x"51c08166",
  3170 => x"87c1fa49",
  3171 => x"c387d1cc",
  3172 => x"d049e0d3",
  3173 => x"e5c08166",
  3174 => x"f949c251",
  3175 => x"ffcb87ef",
  3176 => x"0266d487",
  3177 => x"c387cac0",
  3178 => x"d049e0d3",
  3179 => x"e5c08166",
  3180 => x"d0ffc351",
  3181 => x"c84ac04b",
  3182 => x"fcfc49c0",
  3183 => x"ffc387d4",
  3184 => x"50cb48d7",
  3185 => x"48e0d3c3",
  3186 => x"708066d0",
  3187 => x"bf976e7e",
  3188 => x"c0029949",
  3189 => x"ffc387cc",
  3190 => x"50c548d2",
  3191 => x"976e80c9",
  3192 => x"1ec950bf",
  3193 => x"49d0ffc3",
  3194 => x"c487ccf7",
  3195 => x"f849c086",
  3196 => x"486e87db",
  3197 => x"e7ca50c0",
  3198 => x"0566d487",
  3199 => x"d887f5c2",
  3200 => x"e8c04866",
  3201 => x"c0c105a8",
  3202 => x"4966dc87",
  3203 => x"c0c0c0c1",
  3204 => x"e0c091c0",
  3205 => x"c0d04a66",
  3206 => x"a17292c0",
  3207 => x"9766c449",
  3208 => x"c0c44abf",
  3209 => x"49a17292",
  3210 => x"82c54a6e",
  3211 => x"c04a6a97",
  3212 => x"7248a6e4",
  3213 => x"496e78a1",
  3214 => x"699781c7",
  3215 => x"91c0c449",
  3216 => x"82c84a6e",
  3217 => x"a14a6a97",
  3218 => x"c049744c",
  3219 => x"c08166e4",
  3220 => x"01a966e8",
  3221 => x"c087cbc1",
  3222 => x"c94966e4",
  3223 => x"d01e7131",
  3224 => x"e4fd4966",
  3225 => x"86c487e5",
  3226 => x"8cc14974",
  3227 => x"c0029971",
  3228 => x"66cc87df",
  3229 => x"751ec04d",
  3230 => x"f4defd49",
  3231 => x"751ec187",
  3232 => x"d1ddfd49",
  3233 => x"7486c887",
  3234 => x"718cc149",
  3235 => x"e4ff0599",
  3236 => x"f549c087",
  3237 => x"d3c387f7",
  3238 => x"66d049e0",
  3239 => x"c751c081",
  3240 => x"49c287fe",
  3241 => x"c387e6f5",
  3242 => x"d049e0d3",
  3243 => x"e1c08166",
  3244 => x"87ecc751",
  3245 => x"d4f549c2",
  3246 => x"e0d3c387",
  3247 => x"8166d049",
  3248 => x"c751e5c0",
  3249 => x"66d487da",
  3250 => x"87fdc205",
  3251 => x"c04866d8",
  3252 => x"c105a8ea",
  3253 => x"66dc87c0",
  3254 => x"c0c0c149",
  3255 => x"c091c0c0",
  3256 => x"d04a66e0",
  3257 => x"7292c0c0",
  3258 => x"66c449a1",
  3259 => x"c44abf97",
  3260 => x"a17292c0",
  3261 => x"c54a6e49",
  3262 => x"4a6a9782",
  3263 => x"48a6e4c0",
  3264 => x"6e78a172",
  3265 => x"9781c749",
  3266 => x"c0c44969",
  3267 => x"c84a6e91",
  3268 => x"4a6a9782",
  3269 => x"49744ca1",
  3270 => x"8166e4c0",
  3271 => x"a966e8c0",
  3272 => x"87d3c101",
  3273 => x"c0029c74",
  3274 => x"66cc87fc",
  3275 => x"66e4c04d",
  3276 => x"7131c949",
  3277 => x"fd49751e",
  3278 => x"c387d0e1",
  3279 => x"f249d0ff",
  3280 => x"ffc387eb",
  3281 => x"49751ed0",
  3282 => x"87f4dcfd",
  3283 => x"49751ec1",
  3284 => x"87c2dafd",
  3285 => x"e4c086cc",
  3286 => x"80c14866",
  3287 => x"58a6e8c0",
  3288 => x"ff058cc1",
  3289 => x"49c087c7",
  3290 => x"c387e2f2",
  3291 => x"d049e0d3",
  3292 => x"51c08166",
  3293 => x"c287e9c4",
  3294 => x"87d1f249",
  3295 => x"49e0d3c3",
  3296 => x"c08166d0",
  3297 => x"d7c451e1",
  3298 => x"f149c287",
  3299 => x"d3c387ff",
  3300 => x"66d049e0",
  3301 => x"51e5c081",
  3302 => x"c387c5c4",
  3303 => x"c04bd0ff",
  3304 => x"49c0c84a",
  3305 => x"87eaf4fc",
  3306 => x"48d2ffc3",
  3307 => x"497450c2",
  3308 => x"ffc389c5",
  3309 => x"c35997d8",
  3310 => x"c348ecd2",
  3311 => x"2049d8ff",
  3312 => x"c3412041",
  3313 => x"c348f8d2",
  3314 => x"2049e0ff",
  3315 => x"20412041",
  3316 => x"d0412041",
  3317 => x"f0c04966",
  3318 => x"f2ffc381",
  3319 => x"d3c35997",
  3320 => x"ffc348cc",
  3321 => x"412049f0",
  3322 => x"48d4d3c3",
  3323 => x"49f4ffc3",
  3324 => x"41204120",
  3325 => x"c00266d4",
  3326 => x"ffc387c7",
  3327 => x"ffc148d0",
  3328 => x"c1497450",
  3329 => x"c31e7129",
  3330 => x"ee49d0ff",
  3331 => x"86c487e9",
  3332 => x"f8ef49c0",
  3333 => x"e0d3c387",
  3334 => x"8166d049",
  3335 => x"ffc151c0",
  3336 => x"0566d487",
  3337 => x"c387d2c1",
  3338 => x"c04bd0ff",
  3339 => x"49c0c84a",
  3340 => x"87def2fc",
  3341 => x"48d3ffc3",
  3342 => x"e8c050c8",
  3343 => x"29d04966",
  3344 => x"97d9ffc3",
  3345 => x"66e8c059",
  3346 => x"c329c849",
  3347 => x"5997daff",
  3348 => x"c080c148",
  3349 => x"c25066e8",
  3350 => x"49745080",
  3351 => x"1e7129c1",
  3352 => x"ed49a0f5",
  3353 => x"86c487d1",
  3354 => x"e0ee49c0",
  3355 => x"e0d3c387",
  3356 => x"8166d049",
  3357 => x"e7c051c0",
  3358 => x"e0d3c387",
  3359 => x"8166d049",
  3360 => x"c251e5c0",
  3361 => x"87c5ee49",
  3362 => x"c387d5c0",
  3363 => x"d049e0d3",
  3364 => x"e0c08166",
  3365 => x"ed49c251",
  3366 => x"c3c087f3",
  3367 => x"87c6ee87",
  3368 => x"268ed4ff",
  3369 => x"264c264d",
  3370 => x"004f264b",
  3371 => x"34364354",
  3372 => x"20202020",
  3373 => x"00000000",
  3374 => x"694d6544",
  3375 => x"66695453",
  3376 => x"44482079",
  3377 => x"20302044",
  3378 => x"00000000",
  3379 => x"20323338",
  3380 => x"00000000",
  3381 => x"32313032",
  3382 => x"39323930",
  3383 => x"00000009",
  3384 => x"731e0000",
  3385 => x"ff86e01e",
  3386 => x"c5c848d0",
  3387 => x"48d4ff78",
  3388 => x"1ed078c5",
  3389 => x"494ba6c4",
  3390 => x"87ebf1fc",
  3391 => x"d0ff86c4",
  3392 => x"ca78c448",
  3393 => x"c1496697",
  3394 => x"87c50299",
  3395 => x"e8ec4973",
  3396 => x"268ee087",
  3397 => x"1e4f264b",
  3398 => x"c44ad4ff",
  3399 => x"c448f8d7",
  3400 => x"78bfe4d1",
  3401 => x"ff7affc3",
  3402 => x"78c548d0",
  3403 => x"d1c47ac4",
  3404 => x"4849bfe4",
  3405 => x"7a7028d8",
  3406 => x"28d04871",
  3407 => x"48717a70",
  3408 => x"7a7028c8",
  3409 => x"bfe4d1c4",
  3410 => x"48d0ff7a",
  3411 => x"4f2678c4",
  3412 => x"c44ac01e",
  3413 => x"02bfecd8",
  3414 => x"c44987ca",
  3415 => x"c148ecd8",
  3416 => x"4a1178a1",
  3417 => x"c6059a72",
  3418 => x"ecd8c487",
  3419 => x"7278c048",
  3420 => x"1e4f2648",
  3421 => x"48ecd8c4",
  3422 => x"bfc8f4c3",
  3423 => x"0e4f2678",
  3424 => x"0e5c5b5e",
  3425 => x"d0ff4a71",
  3426 => x"4bd4ff4c",
  3427 => x"d5c17cc5",
  3428 => x"7b66cc7b",
  3429 => x"7cc57cc4",
  3430 => x"c17bd3c1",
  3431 => x"c87cc47b",
  3432 => x"d4c17cc5",
  3433 => x"b749c07b",
  3434 => x"87ca06aa",
  3435 => x"81c17bc0",
  3436 => x"04a9b772",
  3437 => x"7cc487f6",
  3438 => x"d3c17cc5",
  3439 => x"c47bc07b",
  3440 => x"264c267c",
  3441 => x"1e4f264b",
  3442 => x"4b711e73",
  3443 => x"97e0f3c1",
  3444 => x"b7c249bf",
  3445 => x"f3c003a9",
  3446 => x"c41e7387",
  3447 => x"fd49cccc",
  3448 => x"c487d0cb",
  3449 => x"02987086",
  3450 => x"c487e1c0",
  3451 => x"4abfd4cc",
  3452 => x"c0c32aca",
  3453 => x"87ce028a",
  3454 => x"058ac0c1",
  3455 => x"f3c187ce",
  3456 => x"50c048e0",
  3457 => x"f3c187c6",
  3458 => x"50c148e0",
  3459 => x"4f264b26",
  3460 => x"711e731e",
  3461 => x"c6029a4a",
  3462 => x"c4ddc387",
  3463 => x"c378c048",
  3464 => x"49bfc0dd",
  3465 => x"87c0ceff",
  3466 => x"c4029870",
  3467 => x"49d487cd",
  3468 => x"87e8cdff",
  3469 => x"58c4ddc3",
  3470 => x"bfc4ddc3",
  3471 => x"87fbc005",
  3472 => x"49d0d1c4",
  3473 => x"87cedffe",
  3474 => x"04a8b7c0",
  3475 => x"d1c487ce",
  3476 => x"dffe49d0",
  3477 => x"b7c087c0",
  3478 => x"87f203a8",
  3479 => x"bfc4ddc3",
  3480 => x"c4ddc349",
  3481 => x"78a1c148",
  3482 => x"81ccf4c3",
  3483 => x"ddc34811",
  3484 => x"ddc358cc",
  3485 => x"78c048cc",
  3486 => x"c387c0c3",
  3487 => x"02bfccdd",
  3488 => x"c487f5c1",
  3489 => x"fe49d0d1",
  3490 => x"c087cbde",
  3491 => x"cd04a8b7",
  3492 => x"ccddc387",
  3493 => x"88c148bf",
  3494 => x"58d0ddc3",
  3495 => x"d6c487dd",
  3496 => x"ff49bff0",
  3497 => x"7087c1cc",
  3498 => x"cec00298",
  3499 => x"d0d1c487",
  3500 => x"d6dbfe49",
  3501 => x"c4ddc387",
  3502 => x"c378c048",
  3503 => x"05bfc8dd",
  3504 => x"c387f8c1",
  3505 => x"05bfccdd",
  3506 => x"c387f0c1",
  3507 => x"49bfc4dd",
  3508 => x"48c4ddc3",
  3509 => x"c378a1c1",
  3510 => x"1181ccf4",
  3511 => x"c0c2494b",
  3512 => x"ccc00299",
  3513 => x"c1487387",
  3514 => x"ddc398ff",
  3515 => x"cac158d0",
  3516 => x"ccddc387",
  3517 => x"87c3c15b",
  3518 => x"bfc8ddc3",
  3519 => x"87fbc002",
  3520 => x"bfc4ddc3",
  3521 => x"c4ddc349",
  3522 => x"78a1c148",
  3523 => x"81ccf4c3",
  3524 => x"1e496997",
  3525 => x"49d0d1c4",
  3526 => x"87c6dafe",
  3527 => x"ddc386c4",
  3528 => x"c148bfc8",
  3529 => x"ccddc388",
  3530 => x"ccddc358",
  3531 => x"c078c148",
  3532 => x"ff49ecf6",
  3533 => x"c487e5c9",
  3534 => x"2658f4d6",
  3535 => x"004f264b",
  3536 => x"00000000",
  3537 => x"00000000",
  3538 => x"00000000",
  3539 => x"00000000",
  3540 => x"711e731e",
  3541 => x"fbfd494b",
  3542 => x"d1c487f0",
  3543 => x"02bf97f8",
  3544 => x"1ec387cb",
  3545 => x"49c0c0c4",
  3546 => x"c487d4f8",
  3547 => x"fd497386",
  3548 => x"2687d7fb",
  3549 => x"1e4f264b",
  3550 => x"daf61e73",
  3551 => x"49f4c787",
  3552 => x"87d8c8ff",
  3553 => x"ff494b70",
  3554 => x"7087ddc8",
  3555 => x"87cb0598",
  3556 => x"c8ff4973",
  3557 => x"987087d2",
  3558 => x"2687f502",
  3559 => x"0e4f264b",
  3560 => x"5d5c5b5e",
  3561 => x"7186f80e",
  3562 => x"fd4dc04b",
  3563 => x"7087eed4",
  3564 => x"029b734c",
  3565 => x"c187c2c5",
  3566 => x"c148e0f3",
  3567 => x"c41e7350",
  3568 => x"fd49cccc",
  3569 => x"c487ecc3",
  3570 => x"02987086",
  3571 => x"c487ffc3",
  3572 => x"48bfe4d1",
  3573 => x"d1c4b0c1",
  3574 => x"faf458e8",
  3575 => x"d0ffc387",
  3576 => x"ccccc41e",
  3577 => x"c8c9fd49",
  3578 => x"c386c487",
  3579 => x"7ebfdcff",
  3580 => x"c348a6c4",
  3581 => x"78bfe0ff",
  3582 => x"97d0ffc3",
  3583 => x"a9c149bf",
  3584 => x"87cac305",
  3585 => x"bfd4ffc3",
  3586 => x"71b1c149",
  3587 => x"ffcfff48",
  3588 => x"e8d1c498",
  3589 => x"d1ffc358",
  3590 => x"c248bf97",
  3591 => x"c358d0e6",
  3592 => x"49bfd8ff",
  3593 => x"87f2ddfd",
  3594 => x"c0029870",
  3595 => x"ffc387e2",
  3596 => x"ccc41ed0",
  3597 => x"c7fd49cc",
  3598 => x"ffc387f7",
  3599 => x"fd49bfd8",
  3600 => x"c087fbd0",
  3601 => x"e4ffc31e",
  3602 => x"87ccc449",
  3603 => x"4d7086c8",
  3604 => x"d0fd4974",
  3605 => x"1e7387e8",
  3606 => x"49ccccc4",
  3607 => x"87d3c1fd",
  3608 => x"496e86c4",
  3609 => x"87f2dcfd",
  3610 => x"c0029870",
  3611 => x"ffc387e1",
  3612 => x"ccc41ed0",
  3613 => x"c6fd49cc",
  3614 => x"ffc387f7",
  3615 => x"fd49bfdc",
  3616 => x"c087fbcf",
  3617 => x"ffc31ef2",
  3618 => x"cbc349f0",
  3619 => x"7486c887",
  3620 => x"e9cffd49",
  3621 => x"c41e7387",
  3622 => x"fd49cccc",
  3623 => x"c487d4c0",
  3624 => x"fd496686",
  3625 => x"7087f3db",
  3626 => x"e1c00298",
  3627 => x"d0ffc387",
  3628 => x"ccccc41e",
  3629 => x"f8c5fd49",
  3630 => x"e0ffc387",
  3631 => x"cefd49bf",
  3632 => x"f3c087fc",
  3633 => x"fcffc31e",
  3634 => x"87ccc249",
  3635 => x"1ec286c8",
  3636 => x"49c0c0c4",
  3637 => x"c387e8f2",
  3638 => x"c0c0c41e",
  3639 => x"87dff249",
  3640 => x"d1c486c8",
  3641 => x"fe48bfe4",
  3642 => x"e8d1c498",
  3643 => x"87e7f058",
  3644 => x"bfcce6c2",
  3645 => x"d2f5fe49",
  3646 => x"f8487587",
  3647 => x"264d268e",
  3648 => x"264b264c",
  3649 => x"1e731e4f",
  3650 => x"49ca4b71",
  3651 => x"87fedcfc",
  3652 => x"ccc41e73",
  3653 => x"fefc49cc",
  3654 => x"86c487d9",
  3655 => x"c0029870",
  3656 => x"d7c487f0",
  3657 => x"50c148f4",
  3658 => x"bfcce6c2",
  3659 => x"c480c250",
  3660 => x"78bfe4d1",
  3661 => x"50c080db",
  3662 => x"50c080cb",
  3663 => x"50c080cb",
  3664 => x"1ea0c8ff",
  3665 => x"49ccccc4",
  3666 => x"87f4c4fd",
  3667 => x"48c186c4",
  3668 => x"48c087c2",
  3669 => x"4f264b26",
  3670 => x"5c5b5e0e",
  3671 => x"86f40e5d",
  3672 => x"7ec04d71",
  3673 => x"c04866dc",
  3674 => x"a6cc88f0",
  3675 => x"0266dc58",
  3676 => x"7087e6c0",
  3677 => x"f3c10298",
  3678 => x"8cc14c87",
  3679 => x"87ecc102",
  3680 => x"d1c2028c",
  3681 => x"c2028c87",
  3682 => x"8cd087cc",
  3683 => x"87e7c402",
  3684 => x"c4028cc1",
  3685 => x"efc487eb",
  3686 => x"029d7587",
  3687 => x"9787e9c4",
  3688 => x"e3c4026d",
  3689 => x"c41ec287",
  3690 => x"ef49c0c0",
  3691 => x"86c487d1",
  3692 => x"4bc8d8c4",
  3693 => x"49cb4a75",
  3694 => x"87c6dcfc",
  3695 => x"48d3d8c4",
  3696 => x"ccfd50c0",
  3697 => x"d8c487d7",
  3698 => x"d1c458c0",
  3699 => x"c148bfe4",
  3700 => x"e8d1c4b0",
  3701 => x"87ffec58",
  3702 => x"49c8d8c4",
  3703 => x"c487e8ef",
  3704 => x"fd49c8d8",
  3705 => x"c187dee0",
  3706 => x"87dcc37e",
  3707 => x"c01e66c8",
  3708 => x"d7c4ff49",
  3709 => x"4966cc87",
  3710 => x"cc87fcf5",
  3711 => x"49751e66",
  3712 => x"87c8c4ff",
  3713 => x"496686c8",
  3714 => x"c491c8c1",
  3715 => x"c881d0d2",
  3716 => x"c27e6981",
  3717 => x"66c887f2",
  3718 => x"91c8c149",
  3719 => x"48d0d2c4",
  3720 => x"7e708071",
  3721 => x"a680c848",
  3722 => x"4866c458",
  3723 => x"9d7578c0",
  3724 => x"87e6c002",
  3725 => x"cc4c66c8",
  3726 => x"fcd7c494",
  3727 => x"754b7484",
  3728 => x"fc49cb4a",
  3729 => x"cb87fbd9",
  3730 => x"51c049a4",
  3731 => x"66c41e74",
  3732 => x"def9fc49",
  3733 => x"c086c487",
  3734 => x"66c887cb",
  3735 => x"c491cc49",
  3736 => x"c081fcd7",
  3737 => x"f4c9fd51",
  3738 => x"c84a7087",
  3739 => x"91c44966",
  3740 => x"81f8d7c4",
  3741 => x"66c47972",
  3742 => x"dac002bf",
  3743 => x"4966c887",
  3744 => x"c0d089c2",
  3745 => x"70307148",
  3746 => x"e4d1c449",
  3747 => x"b07148bf",
  3748 => x"58e8d1c4",
  3749 => x"c887d9c0",
  3750 => x"89c24966",
  3751 => x"7148c0d0",
  3752 => x"ff497030",
  3753 => x"e4d1c4b9",
  3754 => x"987148bf",
  3755 => x"58e8d1c4",
  3756 => x"7ebf66c4",
  3757 => x"7587d1c0",
  3758 => x"87e3f349",
  3759 => x"c7c07e70",
  3760 => x"f8497587",
  3761 => x"7e7087ff",
  3762 => x"bfe4d1c4",
  3763 => x"c498fe48",
  3764 => x"e958e8d1",
  3765 => x"486e87c1",
  3766 => x"4d268ef4",
  3767 => x"4b264c26",
  3768 => x"731e4f26",
  3769 => x"e4d1c41e",
  3770 => x"c178c148",
  3771 => x"c148e0f3",
  3772 => x"c4c8c150",
  3773 => x"e850c048",
  3774 => x"1ec387dd",
  3775 => x"49c0c0c4",
  3776 => x"c287fce9",
  3777 => x"c0c0c41e",
  3778 => x"87f3e949",
  3779 => x"f4c386c8",
  3780 => x"f249bfe0",
  3781 => x"987087c9",
  3782 => x"87efc105",
  3783 => x"c387f8e7",
  3784 => x"49bfdcf4",
  3785 => x"c387e0ea",
  3786 => x"49bfdcf4",
  3787 => x"87d5dbfd",
  3788 => x"bfe4d1c4",
  3789 => x"c498fe48",
  3790 => x"e758e8d1",
  3791 => x"d0c687d9",
  3792 => x"d7f9fe49",
  3793 => x"494b7087",
  3794 => x"87dcf9fe",
  3795 => x"cc059870",
  3796 => x"fe497387",
  3797 => x"7087d1f9",
  3798 => x"f4ff0298",
  3799 => x"e4d1c487",
  3800 => x"b0c148bf",
  3801 => x"58e8d1c4",
  3802 => x"c187ece6",
  3803 => x"f8fe49e4",
  3804 => x"4b7087ea",
  3805 => x"eff8fe49",
  3806 => x"05987087",
  3807 => x"7387ccc0",
  3808 => x"e3f8fe49",
  3809 => x"02987087",
  3810 => x"c487f4ff",
  3811 => x"48bfe4d1",
  3812 => x"d1c498fe",
  3813 => x"fee558e8",
  3814 => x"fbcfff87",
  3815 => x"dac7fe87",
  3816 => x"e949c187",
  3817 => x"48c087ea",
  3818 => x"4f264b26",
  3819 => x"711e731e",
  3820 => x"cfc4ff4b",
  3821 => x"fe497387",
  3822 => x"2687d0cf",
  3823 => x"0e4f264b",
  3824 => x"0e5c5b5e",
  3825 => x"ffc186fc",
  3826 => x"4b6e4cff",
  3827 => x"ffe849c0",
  3828 => x"deedfe87",
  3829 => x"dcf9fe87",
  3830 => x"87c6e487",
  3831 => x"99744973",
  3832 => x"997183c1",
  3833 => x"fd87e505",
  3834 => x"7087f9ff",
  3835 => x"eed4fe49",
  3836 => x"87d8ff87",
  3837 => x"4c268efc",
  3838 => x"4f264b26",
  3839 => x"f5f2ebf4",
  3840 => x"0c040605",
  3841 => x"0a830b03",
  3842 => x"00000066",
  3843 => x"00da005a",
  3844 => x"08948000",
  3845 => x"00788005",
  3846 => x"00018002",
  3847 => x"00098003",
  3848 => x"00008004",
  3849 => x"08918001",
  3850 => x"00000026",
  3851 => x"0000001d",
  3852 => x"0000001c",
  3853 => x"00000025",
  3854 => x"0000001a",
  3855 => x"0000001b",
  3856 => x"00000024",
  3857 => x"00000112",
  3858 => x"0000002e",
  3859 => x"0000002d",
  3860 => x"00000023",
  3861 => x"00000036",
  3862 => x"00000021",
  3863 => x"0000002b",
  3864 => x"0000002c",
  3865 => x"00000022",
  3866 => x"006c003d",
  3867 => x"00000035",
  3868 => x"00000034",
  3869 => x"0075003e",
  3870 => x"00000032",
  3871 => x"00000033",
  3872 => x"006b003c",
  3873 => x"0000002a",
  3874 => x"007d0046",
  3875 => x"00730043",
  3876 => x"0069003b",
  3877 => x"00ca0045",
  3878 => x"0070003a",
  3879 => x"00720042",
  3880 => x"00740044",
  3881 => x"00000031",
  3882 => x"00000055",
  3883 => x"007c004d",
  3884 => x"007a004b",
  3885 => x"0000007b",
  3886 => x"00710049",
  3887 => x"0084004c",
  3888 => x"00770054",
  3889 => x"00000041",
  3890 => x"00000061",
  3891 => x"007c005b",
  3892 => x"00000052",
  3893 => x"000000f1",
  3894 => x"00000259",
  3895 => x"005d000e",
  3896 => x"0000005d",
  3897 => x"0079004a",
  3898 => x"00000016",
  3899 => x"00070076",
  3900 => x"000d0414",
  3901 => x"0000001e",
  3902 => x"00000029",
  3903 => x"00000011",
  3904 => x"00000015",
  3905 => x"00004000",
  3906 => x"00003d24",
  3907 => x"0882ff01",
  3908 => x"64f3c8f3",
  3909 => x"01f250f3",
  3910 => x"00f40181",
  3911 => x"00003f90",
  3912 => x"00003f9c",
  3913 => x"72617441",
  3914 => x"54532069",
  3915 => x"31503b3b",
  3916 => x"6f74532c",
  3917 => x"65676172",
  3918 => x"5331503b",
  3919 => x"532c5530",
  3920 => x"462c2054",
  3921 => x"70706f6c",
  3922 => x"3a412079",
  3923 => x"5331503b",
  3924 => x"532c5531",
  3925 => x"462c2054",
  3926 => x"70706f6c",
  3927 => x"3a422079",
  3928 => x"4f31503b",
  3929 => x"572c3736",
  3930 => x"65746972",
  3931 => x"6f727020",
  3932 => x"74636574",
  3933 => x"66664f2c",
  3934 => x"2c3a412c",
  3935 => x"422c3a42",
  3936 => x"3b68746f",
  3937 => x"414f3150",
  3938 => x"61482c42",
  3939 => x"64206472",
  3940 => x"736b7369",
  3941 => x"6e6f4e2c",
  3942 => x"6e552c65",
  3943 => x"30207469",
  3944 => x"696e552c",
  3945 => x"2c312074",
  3946 => x"68746f42",
  3947 => x"5331503b",
  3948 => x"482c5532",
  3949 => x"48564644",
  3950 => x"61482c44",
  3951 => x"69666472",
  3952 => x"3020656c",
  3953 => x"5331503b",
  3954 => x"482c5533",
  3955 => x"48564644",
  3956 => x"61482c44",
  3957 => x"69666472",
  3958 => x"3120656c",
  3959 => x"2c32503b",
  3960 => x"74737953",
  3961 => x"503b6d65",
  3962 => x"4f4e4f32",
  3963 => x"6968432c",
  3964 => x"74657370",
  3965 => x"2c54532c",
  3966 => x"2c455453",
  3967 => x"6167654d",
  3968 => x"2c455453",
  3969 => x"72455453",
  3970 => x"7364696f",
  3971 => x"4f32503b",
  3972 => x"54532c4a",
  3973 => x"696c4220",
  3974 => x"72657474",
  3975 => x"66664f2c",
  3976 => x"3b6e4f2c",
  3977 => x"314f3250",
  3978 => x"41522c33",
  3979 => x"6e28204d",
  3980 => x"20646565",
  3981 => x"64726148",
  3982 => x"73655220",
  3983 => x"2c297465",
  3984 => x"4b323135",
  3985 => x"424d312c",
  3986 => x"424d322c",
  3987 => x"424d342c",
  3988 => x"424d382c",
  3989 => x"4d34312c",
  3990 => x"32503b42",
  3991 => x"4d492c46",
  3992 => x"4d4f5247",
  3993 => x"616f4c2c",
  3994 => x"4f522064",
  3995 => x"32503b4d",
  3996 => x"49422c46",
  3997 => x"4354534e",
  3998 => x"616f4c2c",
  3999 => x"61432064",
  4000 => x"69727472",
  4001 => x"3b656764",
  4002 => x"532c3350",
  4003 => x"646e756f",
  4004 => x"56202620",
  4005 => x"6f656469",
  4006 => x"4f33503b",
  4007 => x"69562c38",
  4008 => x"206f6564",
  4009 => x"65646f6d",
  4010 => x"6e6f4d2c",
  4011 => x"6f432c6f",
  4012 => x"72756f6c",
  4013 => x"4f33503b",
  4014 => x"69562c53",
  4015 => x"676e696b",
  4016 => x"314d532f",
  4017 => x"4f2c3439",
  4018 => x"4f2c6666",
  4019 => x"33503b6e",
  4020 => x"2c4c4b4f",
  4021 => x"6e616353",
  4022 => x"656e696c",
  4023 => x"664f2c73",
  4024 => x"35322c66",
  4025 => x"30352c25",
  4026 => x"35372c25",
  4027 => x"33503b25",
  4028 => x"432c544f",
  4029 => x"6f706d6f",
  4030 => x"65746973",
  4031 => x"656c6220",
  4032 => x"4f2c646e",
  4033 => x"4f2c6666",
  4034 => x"33503b6e",
  4035 => x"532c4d4f",
  4036 => x"65726574",
  4037 => x"6f73206f",
  4038 => x"2c646e75",
  4039 => x"2c66664f",
  4040 => x"503b6e4f",
  4041 => x"2c554f33",
  4042 => x"69657453",
  4043 => x"7265626e",
  4044 => x"6f642067",
  4045 => x"656c676e",
  4046 => x"66664f2c",
  4047 => x"3b6e4f2c",
  4048 => x"432c4353",
  4049 => x"4c2c4746",
  4050 => x"2064616f",
  4051 => x"666e6f63",
  4052 => x"533b6769",
  4053 => x"46432c44",
  4054 => x"61532c47",
  4055 => x"63206576",
  4056 => x"69666e6f",
  4057 => x"30543b67",
  4058 => x"7365522c",
  4059 => x"28207465",
  4060 => x"646c6f48",
  4061 => x"726f6620",
  4062 => x"72616820",
  4063 => x"65722064",
  4064 => x"29746573",
  4065 => x"762c563b",
  4066 => x"30342e33",
  4067 => x"0000002e",
  4068 => x"20534f54",
  4069 => x"20202020",
  4070 => x"00474d49",
  4071 => x"5453494d",
  4072 => x"20595245",
  4073 => x"00474643",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
