
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"d8",x"c4",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f0",x"d8",x"c4"),
    14 => (x"48",x"e8",x"fe",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fc",x"f1"),
    19 => (x"fc",x"1e",x"87",x"fd"),
    20 => (x"ff",x"4a",x"71",x"86"),
    21 => (x"48",x"69",x"49",x"c0"),
    22 => (x"70",x"98",x"c0",x"c4"),
    23 => (x"02",x"98",x"48",x"7e"),
    24 => (x"79",x"72",x"87",x"f4"),
    25 => (x"26",x"8e",x"fc",x"48"),
    26 => (x"1e",x"72",x"1e",x"4f"),
    27 => (x"48",x"12",x"1e",x"73"),
    28 => (x"87",x"ca",x"02",x"11"),
    29 => (x"98",x"df",x"c3",x"4b"),
    30 => (x"02",x"88",x"73",x"9b"),
    31 => (x"4b",x"26",x"87",x"f0"),
    32 => (x"4f",x"26",x"4a",x"26"),
    33 => (x"72",x"1e",x"73",x"1e"),
    34 => (x"04",x"8b",x"c1",x"1e"),
    35 => (x"48",x"12",x"87",x"ca"),
    36 => (x"87",x"c4",x"02",x"11"),
    37 => (x"87",x"f1",x"02",x"88"),
    38 => (x"4b",x"26",x"4a",x"26"),
    39 => (x"74",x"1e",x"4f",x"26"),
    40 => (x"72",x"1e",x"73",x"1e"),
    41 => (x"04",x"8b",x"c1",x"1e"),
    42 => (x"48",x"12",x"87",x"d0"),
    43 => (x"87",x"ca",x"02",x"11"),
    44 => (x"98",x"df",x"c3",x"4c"),
    45 => (x"02",x"88",x"74",x"9c"),
    46 => (x"4a",x"26",x"87",x"eb"),
    47 => (x"4c",x"26",x"4b",x"26"),
    48 => (x"73",x"1e",x"4f",x"26"),
    49 => (x"a9",x"73",x"81",x"48"),
    50 => (x"12",x"87",x"c5",x"02"),
    51 => (x"87",x"f6",x"05",x"53"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"a9",x"73",x"81",x"48"),
    54 => (x"f9",x"53",x"72",x"05"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"9a",x"72",x"1e",x"73"),
    57 => (x"87",x"e7",x"c0",x"02"),
    58 => (x"4b",x"c1",x"48",x"c0"),
    59 => (x"d1",x"06",x"a9",x"72"),
    60 => (x"06",x"82",x"72",x"87"),
    61 => (x"83",x"73",x"87",x"c9"),
    62 => (x"f4",x"01",x"a9",x"72"),
    63 => (x"c1",x"87",x"c3",x"87"),
    64 => (x"a9",x"72",x"3a",x"b2"),
    65 => (x"80",x"73",x"89",x"03"),
    66 => (x"2b",x"2a",x"c1",x"07"),
    67 => (x"26",x"87",x"f3",x"05"),
    68 => (x"1e",x"4f",x"26",x"4b"),
    69 => (x"4d",x"c4",x"1e",x"75"),
    70 => (x"04",x"a1",x"b7",x"71"),
    71 => (x"81",x"c1",x"b9",x"ff"),
    72 => (x"72",x"07",x"bd",x"c3"),
    73 => (x"ff",x"04",x"a2",x"b7"),
    74 => (x"c1",x"82",x"c1",x"ba"),
    75 => (x"ee",x"fe",x"07",x"bd"),
    76 => (x"04",x"2d",x"c1",x"87"),
    77 => (x"80",x"c1",x"b8",x"ff"),
    78 => (x"ff",x"04",x"2d",x"07"),
    79 => (x"07",x"81",x"c1",x"b9"),
    80 => (x"4f",x"26",x"4d",x"26"),
    81 => (x"71",x"1e",x"73",x"1e"),
    82 => (x"4b",x"66",x"c8",x"4a"),
    83 => (x"71",x"8b",x"c1",x"49"),
    84 => (x"87",x"cf",x"02",x"99"),
    85 => (x"d4",x"ff",x"48",x"12"),
    86 => (x"49",x"73",x"78",x"08"),
    87 => (x"99",x"71",x"8b",x"c1"),
    88 => (x"26",x"87",x"f1",x"05"),
    89 => (x"0e",x"4f",x"26",x"4b"),
    90 => (x"0e",x"5c",x"5b",x"5e"),
    91 => (x"d4",x"ff",x"4a",x"71"),
    92 => (x"4b",x"66",x"cc",x"4c"),
    93 => (x"71",x"8b",x"c1",x"49"),
    94 => (x"87",x"ce",x"02",x"99"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"c1",x"49",x"73",x"52"),
    97 => (x"05",x"99",x"71",x"8b"),
    98 => (x"4c",x"26",x"87",x"f2"),
    99 => (x"4f",x"26",x"4b",x"26"),
   100 => (x"ff",x"1e",x"73",x"1e"),
   101 => (x"ff",x"c3",x"4b",x"d4"),
   102 => (x"c3",x"4a",x"6b",x"7b"),
   103 => (x"49",x"6b",x"7b",x"ff"),
   104 => (x"b1",x"72",x"32",x"c8"),
   105 => (x"6b",x"7b",x"ff",x"c3"),
   106 => (x"71",x"31",x"c8",x"4a"),
   107 => (x"7b",x"ff",x"c3",x"b2"),
   108 => (x"32",x"c8",x"49",x"6b"),
   109 => (x"48",x"71",x"b1",x"72"),
   110 => (x"4f",x"26",x"4b",x"26"),
   111 => (x"5c",x"5b",x"5e",x"0e"),
   112 => (x"4d",x"71",x"0e",x"5d"),
   113 => (x"75",x"4c",x"d4",x"ff"),
   114 => (x"98",x"ff",x"c3",x"48"),
   115 => (x"fe",x"c3",x"7c",x"70"),
   116 => (x"c8",x"05",x"bf",x"e8"),
   117 => (x"48",x"66",x"d0",x"87"),
   118 => (x"a6",x"d4",x"30",x"c9"),
   119 => (x"49",x"66",x"d0",x"58"),
   120 => (x"48",x"71",x"29",x"d8"),
   121 => (x"70",x"98",x"ff",x"c3"),
   122 => (x"49",x"66",x"d0",x"7c"),
   123 => (x"48",x"71",x"29",x"d0"),
   124 => (x"70",x"98",x"ff",x"c3"),
   125 => (x"49",x"66",x"d0",x"7c"),
   126 => (x"48",x"71",x"29",x"c8"),
   127 => (x"70",x"98",x"ff",x"c3"),
   128 => (x"48",x"66",x"d0",x"7c"),
   129 => (x"70",x"98",x"ff",x"c3"),
   130 => (x"d0",x"49",x"75",x"7c"),
   131 => (x"c3",x"48",x"71",x"29"),
   132 => (x"7c",x"70",x"98",x"ff"),
   133 => (x"f0",x"c9",x"4b",x"6c"),
   134 => (x"ff",x"c3",x"4a",x"ff"),
   135 => (x"87",x"cf",x"05",x"ab"),
   136 => (x"6c",x"7c",x"71",x"49"),
   137 => (x"02",x"8a",x"c1",x"4b"),
   138 => (x"ab",x"71",x"87",x"c5"),
   139 => (x"73",x"87",x"f2",x"02"),
   140 => (x"26",x"4d",x"26",x"48"),
   141 => (x"26",x"4b",x"26",x"4c"),
   142 => (x"49",x"c0",x"1e",x"4f"),
   143 => (x"c3",x"48",x"d4",x"ff"),
   144 => (x"81",x"c1",x"78",x"ff"),
   145 => (x"a9",x"b7",x"c8",x"c3"),
   146 => (x"26",x"87",x"f1",x"04"),
   147 => (x"5b",x"5e",x"0e",x"4f"),
   148 => (x"c0",x"0e",x"5d",x"5c"),
   149 => (x"f7",x"c1",x"f0",x"ff"),
   150 => (x"c0",x"c0",x"c1",x"4d"),
   151 => (x"4b",x"c0",x"c0",x"c0"),
   152 => (x"c4",x"87",x"d6",x"ff"),
   153 => (x"c0",x"4c",x"df",x"f8"),
   154 => (x"fd",x"49",x"75",x"1e"),
   155 => (x"86",x"c4",x"87",x"ce"),
   156 => (x"c0",x"05",x"a8",x"c1"),
   157 => (x"d4",x"ff",x"87",x"e5"),
   158 => (x"78",x"ff",x"c3",x"48"),
   159 => (x"e1",x"c0",x"1e",x"73"),
   160 => (x"49",x"e9",x"c1",x"f0"),
   161 => (x"c4",x"87",x"f5",x"fc"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"d4",x"ff",x"87",x"ca"),
   164 => (x"78",x"ff",x"c3",x"48"),
   165 => (x"87",x"cb",x"48",x"c1"),
   166 => (x"c1",x"87",x"de",x"fe"),
   167 => (x"c6",x"ff",x"05",x"8c"),
   168 => (x"26",x"48",x"c0",x"87"),
   169 => (x"26",x"4c",x"26",x"4d"),
   170 => (x"0e",x"4f",x"26",x"4b"),
   171 => (x"0e",x"5c",x"5b",x"5e"),
   172 => (x"c1",x"f0",x"ff",x"c0"),
   173 => (x"d4",x"ff",x"4c",x"c1"),
   174 => (x"78",x"ff",x"c3",x"48"),
   175 => (x"1e",x"c0",x"4b",x"d3"),
   176 => (x"f7",x"fb",x"49",x"74"),
   177 => (x"70",x"86",x"c4",x"87"),
   178 => (x"87",x"ca",x"05",x"98"),
   179 => (x"c3",x"48",x"d4",x"ff"),
   180 => (x"48",x"c1",x"78",x"ff"),
   181 => (x"e0",x"fd",x"87",x"ca"),
   182 => (x"05",x"8b",x"c1",x"87"),
   183 => (x"48",x"c0",x"87",x"e0"),
   184 => (x"4b",x"26",x"4c",x"26"),
   185 => (x"5e",x"0e",x"4f",x"26"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"c4",x"fd",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"fb",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"e0",x"fe"),
   195 => (x"87",x"e2",x"c1",x"48"),
   196 => (x"70",x"87",x"fd",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fe",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"c9"),
   201 => (x"75",x"87",x"cb",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"de",x"fc"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"fc",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"d5",x"48",x"c1",x"87"),
   215 => (x"d1",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"48",x"c0",x"87",x"c4"),
   218 => (x"8c",x"c1",x"87",x"c8"),
   219 => (x"87",x"fc",x"fe",x"05"),
   220 => (x"4d",x"26",x"48",x"c0"),
   221 => (x"4b",x"26",x"4c",x"26"),
   222 => (x"5e",x"0e",x"4f",x"26"),
   223 => (x"0e",x"5d",x"5c",x"5b"),
   224 => (x"c0",x"4d",x"d0",x"ff"),
   225 => (x"c0",x"c1",x"d0",x"e5"),
   226 => (x"e8",x"fe",x"c3",x"4c"),
   227 => (x"c7",x"78",x"c1",x"48"),
   228 => (x"fa",x"7d",x"c2",x"4b"),
   229 => (x"7d",x"c3",x"87",x"e3"),
   230 => (x"49",x"74",x"1e",x"c0"),
   231 => (x"c4",x"87",x"dd",x"f8"),
   232 => (x"05",x"a8",x"c1",x"86"),
   233 => (x"c2",x"4b",x"87",x"c1"),
   234 => (x"87",x"c5",x"05",x"ab"),
   235 => (x"f6",x"c0",x"48",x"c0"),
   236 => (x"05",x"8b",x"c1",x"87"),
   237 => (x"fc",x"87",x"da",x"ff"),
   238 => (x"fe",x"c3",x"87",x"ec"),
   239 => (x"98",x"70",x"58",x"ec"),
   240 => (x"c1",x"87",x"cd",x"05"),
   241 => (x"f0",x"ff",x"c0",x"1e"),
   242 => (x"f7",x"49",x"d0",x"c1"),
   243 => (x"86",x"c4",x"87",x"ee"),
   244 => (x"c3",x"48",x"d4",x"ff"),
   245 => (x"e8",x"c4",x"78",x"ff"),
   246 => (x"f0",x"fe",x"c3",x"87"),
   247 => (x"ff",x"7d",x"c2",x"58"),
   248 => (x"ff",x"c3",x"48",x"d4"),
   249 => (x"26",x"48",x"c1",x"78"),
   250 => (x"26",x"4c",x"26",x"4d"),
   251 => (x"0e",x"4f",x"26",x"4b"),
   252 => (x"5d",x"5c",x"5b",x"5e"),
   253 => (x"c3",x"4d",x"71",x"0e"),
   254 => (x"d4",x"ff",x"4c",x"ff"),
   255 => (x"ff",x"7b",x"74",x"4b"),
   256 => (x"c3",x"c4",x"48",x"d0"),
   257 => (x"75",x"7b",x"74",x"78"),
   258 => (x"f0",x"ff",x"c0",x"1e"),
   259 => (x"f6",x"49",x"d8",x"c1"),
   260 => (x"86",x"c4",x"87",x"ea"),
   261 => (x"c5",x"02",x"98",x"70"),
   262 => (x"c0",x"48",x"c1",x"87"),
   263 => (x"7b",x"74",x"87",x"ee"),
   264 => (x"c8",x"7b",x"fe",x"c3"),
   265 => (x"66",x"d4",x"1e",x"c0"),
   266 => (x"87",x"d8",x"f4",x"49"),
   267 => (x"7b",x"74",x"86",x"c4"),
   268 => (x"7b",x"74",x"7b",x"74"),
   269 => (x"4a",x"e0",x"da",x"d8"),
   270 => (x"05",x"6b",x"7b",x"74"),
   271 => (x"8a",x"c1",x"87",x"c5"),
   272 => (x"74",x"87",x"f5",x"05"),
   273 => (x"48",x"d0",x"ff",x"7b"),
   274 => (x"48",x"c0",x"78",x"c2"),
   275 => (x"4c",x"26",x"4d",x"26"),
   276 => (x"4f",x"26",x"4b",x"26"),
   277 => (x"5c",x"5b",x"5e",x"0e"),
   278 => (x"86",x"fc",x"0e",x"5d"),
   279 => (x"d4",x"ff",x"4b",x"71"),
   280 => (x"c5",x"7e",x"c0",x"4c"),
   281 => (x"4a",x"df",x"cd",x"ee"),
   282 => (x"6c",x"7c",x"ff",x"c3"),
   283 => (x"a8",x"fe",x"c3",x"48"),
   284 => (x"87",x"f8",x"c0",x"05"),
   285 => (x"9b",x"73",x"4d",x"74"),
   286 => (x"d4",x"87",x"cc",x"02"),
   287 => (x"49",x"73",x"1e",x"66"),
   288 => (x"c4",x"87",x"e4",x"f3"),
   289 => (x"ff",x"87",x"d4",x"86"),
   290 => (x"d1",x"c4",x"48",x"d0"),
   291 => (x"4a",x"66",x"d4",x"78"),
   292 => (x"c1",x"7d",x"ff",x"c3"),
   293 => (x"87",x"f8",x"05",x"8a"),
   294 => (x"c3",x"5a",x"a6",x"d8"),
   295 => (x"73",x"7c",x"7c",x"ff"),
   296 => (x"87",x"c5",x"05",x"9b"),
   297 => (x"d0",x"48",x"d0",x"ff"),
   298 => (x"7e",x"4a",x"c1",x"78"),
   299 => (x"fe",x"05",x"8a",x"c1"),
   300 => (x"48",x"6e",x"87",x"f6"),
   301 => (x"4d",x"26",x"8e",x"fc"),
   302 => (x"4b",x"26",x"4c",x"26"),
   303 => (x"73",x"1e",x"4f",x"26"),
   304 => (x"c0",x"4a",x"71",x"1e"),
   305 => (x"48",x"d4",x"ff",x"4b"),
   306 => (x"ff",x"78",x"ff",x"c3"),
   307 => (x"c3",x"c4",x"48",x"d0"),
   308 => (x"48",x"d4",x"ff",x"78"),
   309 => (x"72",x"78",x"ff",x"c3"),
   310 => (x"f0",x"ff",x"c0",x"1e"),
   311 => (x"f3",x"49",x"d1",x"c1"),
   312 => (x"86",x"c4",x"87",x"da"),
   313 => (x"d2",x"05",x"98",x"70"),
   314 => (x"1e",x"c0",x"c8",x"87"),
   315 => (x"fd",x"49",x"66",x"cc"),
   316 => (x"86",x"c4",x"87",x"e2"),
   317 => (x"d0",x"ff",x"4b",x"70"),
   318 => (x"73",x"78",x"c2",x"48"),
   319 => (x"26",x"4b",x"26",x"48"),
   320 => (x"5b",x"5e",x"0e",x"4f"),
   321 => (x"c0",x"0e",x"5d",x"5c"),
   322 => (x"f0",x"ff",x"c0",x"1e"),
   323 => (x"f2",x"49",x"c9",x"c1"),
   324 => (x"1e",x"d2",x"87",x"ea"),
   325 => (x"49",x"f0",x"fe",x"c3"),
   326 => (x"c8",x"87",x"f9",x"fc"),
   327 => (x"c1",x"4c",x"c0",x"86"),
   328 => (x"ac",x"b7",x"d2",x"84"),
   329 => (x"c3",x"87",x"f8",x"04"),
   330 => (x"bf",x"97",x"f0",x"fe"),
   331 => (x"99",x"c0",x"c3",x"49"),
   332 => (x"05",x"a9",x"c0",x"c1"),
   333 => (x"c3",x"87",x"e7",x"c0"),
   334 => (x"bf",x"97",x"f7",x"fe"),
   335 => (x"c3",x"31",x"d0",x"49"),
   336 => (x"bf",x"97",x"f8",x"fe"),
   337 => (x"72",x"32",x"c8",x"4a"),
   338 => (x"f9",x"fe",x"c3",x"b1"),
   339 => (x"b1",x"4a",x"bf",x"97"),
   340 => (x"ff",x"cf",x"4c",x"71"),
   341 => (x"c1",x"9c",x"ff",x"ff"),
   342 => (x"c1",x"34",x"ca",x"84"),
   343 => (x"fe",x"c3",x"87",x"e7"),
   344 => (x"49",x"bf",x"97",x"f9"),
   345 => (x"99",x"c6",x"31",x"c1"),
   346 => (x"97",x"fa",x"fe",x"c3"),
   347 => (x"b7",x"c7",x"4a",x"bf"),
   348 => (x"c3",x"b1",x"72",x"2a"),
   349 => (x"bf",x"97",x"f5",x"fe"),
   350 => (x"9d",x"cf",x"4d",x"4a"),
   351 => (x"97",x"f6",x"fe",x"c3"),
   352 => (x"9a",x"c3",x"4a",x"bf"),
   353 => (x"fe",x"c3",x"32",x"ca"),
   354 => (x"4b",x"bf",x"97",x"f7"),
   355 => (x"b2",x"73",x"33",x"c2"),
   356 => (x"97",x"f8",x"fe",x"c3"),
   357 => (x"c0",x"c3",x"4b",x"bf"),
   358 => (x"2b",x"b7",x"c6",x"9b"),
   359 => (x"81",x"c2",x"b2",x"73"),
   360 => (x"30",x"71",x"48",x"c1"),
   361 => (x"48",x"c1",x"49",x"70"),
   362 => (x"4d",x"70",x"30",x"75"),
   363 => (x"84",x"c1",x"4c",x"72"),
   364 => (x"c0",x"c8",x"94",x"71"),
   365 => (x"cc",x"06",x"ad",x"b7"),
   366 => (x"b7",x"34",x"c1",x"87"),
   367 => (x"b7",x"c0",x"c8",x"2d"),
   368 => (x"f4",x"ff",x"01",x"ad"),
   369 => (x"26",x"48",x"74",x"87"),
   370 => (x"26",x"4c",x"26",x"4d"),
   371 => (x"0e",x"4f",x"26",x"4b"),
   372 => (x"5d",x"5c",x"5b",x"5e"),
   373 => (x"c4",x"86",x"f8",x"0e"),
   374 => (x"c0",x"48",x"d8",x"c7"),
   375 => (x"d0",x"ff",x"c3",x"78"),
   376 => (x"fb",x"49",x"c0",x"1e"),
   377 => (x"86",x"c4",x"87",x"d8"),
   378 => (x"c5",x"05",x"98",x"70"),
   379 => (x"c9",x"48",x"c0",x"87"),
   380 => (x"4d",x"c0",x"87",x"c0"),
   381 => (x"c2",x"c1",x"7e",x"c1"),
   382 => (x"c4",x"49",x"bf",x"d0"),
   383 => (x"71",x"4a",x"c6",x"c0"),
   384 => (x"ff",x"e9",x"4b",x"c8"),
   385 => (x"05",x"98",x"70",x"87"),
   386 => (x"7e",x"c0",x"87",x"c2"),
   387 => (x"bf",x"cc",x"c2",x"c1"),
   388 => (x"e2",x"c0",x"c4",x"49"),
   389 => (x"4b",x"c8",x"71",x"4a"),
   390 => (x"70",x"87",x"e9",x"e9"),
   391 => (x"87",x"c2",x"05",x"98"),
   392 => (x"02",x"6e",x"7e",x"c0"),
   393 => (x"c4",x"87",x"fd",x"c0"),
   394 => (x"4d",x"bf",x"d6",x"c6"),
   395 => (x"9f",x"ce",x"c7",x"c4"),
   396 => (x"c5",x"48",x"7e",x"bf"),
   397 => (x"05",x"a8",x"ea",x"d6"),
   398 => (x"c6",x"c4",x"87",x"c7"),
   399 => (x"ce",x"4d",x"bf",x"d6"),
   400 => (x"ca",x"48",x"6e",x"87"),
   401 => (x"02",x"a8",x"d5",x"e9"),
   402 => (x"48",x"c0",x"87",x"c5"),
   403 => (x"c3",x"87",x"e3",x"c7"),
   404 => (x"75",x"1e",x"d0",x"ff"),
   405 => (x"87",x"e6",x"f9",x"49"),
   406 => (x"98",x"70",x"86",x"c4"),
   407 => (x"c0",x"87",x"c5",x"05"),
   408 => (x"87",x"ce",x"c7",x"48"),
   409 => (x"bf",x"cc",x"c2",x"c1"),
   410 => (x"e2",x"c0",x"c4",x"49"),
   411 => (x"4b",x"c8",x"71",x"4a"),
   412 => (x"70",x"87",x"d1",x"e8"),
   413 => (x"87",x"c8",x"05",x"98"),
   414 => (x"48",x"d8",x"c7",x"c4"),
   415 => (x"87",x"da",x"78",x"c1"),
   416 => (x"bf",x"d0",x"c2",x"c1"),
   417 => (x"c6",x"c0",x"c4",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"f5",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c6",x"48",x"c0",x"87"),
   422 => (x"c7",x"c4",x"87",x"d8"),
   423 => (x"49",x"bf",x"97",x"ce"),
   424 => (x"05",x"a9",x"d5",x"c1"),
   425 => (x"c4",x"87",x"cd",x"c0"),
   426 => (x"bf",x"97",x"cf",x"c7"),
   427 => (x"a9",x"ea",x"c2",x"49"),
   428 => (x"87",x"c5",x"c0",x"02"),
   429 => (x"f9",x"c5",x"48",x"c0"),
   430 => (x"d0",x"ff",x"c3",x"87"),
   431 => (x"48",x"7e",x"bf",x"97"),
   432 => (x"02",x"a8",x"e9",x"c3"),
   433 => (x"6e",x"87",x"ce",x"c0"),
   434 => (x"a8",x"eb",x"c3",x"48"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dd",x"c5",x"48",x"c0"),
   437 => (x"db",x"ff",x"c3",x"87"),
   438 => (x"99",x"49",x"bf",x"97"),
   439 => (x"87",x"cc",x"c0",x"05"),
   440 => (x"97",x"dc",x"ff",x"c3"),
   441 => (x"a9",x"c2",x"49",x"bf"),
   442 => (x"87",x"c5",x"c0",x"02"),
   443 => (x"c1",x"c5",x"48",x"c0"),
   444 => (x"dd",x"ff",x"c3",x"87"),
   445 => (x"c4",x"48",x"bf",x"97"),
   446 => (x"70",x"58",x"d4",x"c7"),
   447 => (x"88",x"c1",x"48",x"4c"),
   448 => (x"58",x"d8",x"c7",x"c4"),
   449 => (x"97",x"de",x"ff",x"c3"),
   450 => (x"81",x"75",x"49",x"bf"),
   451 => (x"97",x"df",x"ff",x"c3"),
   452 => (x"32",x"c8",x"4a",x"bf"),
   453 => (x"c4",x"7e",x"a1",x"72"),
   454 => (x"6e",x"48",x"e8",x"cb"),
   455 => (x"e0",x"ff",x"c3",x"78"),
   456 => (x"c8",x"48",x"bf",x"97"),
   457 => (x"c7",x"c4",x"58",x"a6"),
   458 => (x"c2",x"02",x"bf",x"d8"),
   459 => (x"c2",x"c1",x"87",x"cf"),
   460 => (x"c4",x"49",x"bf",x"cc"),
   461 => (x"71",x"4a",x"e2",x"c0"),
   462 => (x"c7",x"e5",x"4b",x"c8"),
   463 => (x"02",x"98",x"70",x"87"),
   464 => (x"c0",x"87",x"c5",x"c0"),
   465 => (x"87",x"ea",x"c3",x"48"),
   466 => (x"bf",x"d0",x"c7",x"c4"),
   467 => (x"fc",x"cb",x"c4",x"4c"),
   468 => (x"f5",x"ff",x"c3",x"5c"),
   469 => (x"c8",x"49",x"bf",x"97"),
   470 => (x"f4",x"ff",x"c3",x"31"),
   471 => (x"a1",x"4a",x"bf",x"97"),
   472 => (x"f6",x"ff",x"c3",x"49"),
   473 => (x"d0",x"4a",x"bf",x"97"),
   474 => (x"49",x"a1",x"72",x"32"),
   475 => (x"97",x"f7",x"ff",x"c3"),
   476 => (x"32",x"d8",x"4a",x"bf"),
   477 => (x"c4",x"49",x"a1",x"72"),
   478 => (x"cb",x"c4",x"91",x"66"),
   479 => (x"c4",x"81",x"bf",x"e8"),
   480 => (x"c3",x"59",x"f0",x"cb"),
   481 => (x"bf",x"97",x"fd",x"ff"),
   482 => (x"c3",x"32",x"c8",x"4a"),
   483 => (x"bf",x"97",x"fc",x"ff"),
   484 => (x"c3",x"4a",x"a2",x"4b"),
   485 => (x"bf",x"97",x"fe",x"ff"),
   486 => (x"73",x"33",x"d0",x"4b"),
   487 => (x"ff",x"c3",x"4a",x"a2"),
   488 => (x"4b",x"bf",x"97",x"ff"),
   489 => (x"33",x"d8",x"9b",x"cf"),
   490 => (x"c4",x"4a",x"a2",x"73"),
   491 => (x"c2",x"5a",x"f4",x"cb"),
   492 => (x"c4",x"92",x"74",x"8a"),
   493 => (x"72",x"48",x"f4",x"cb"),
   494 => (x"c1",x"c1",x"78",x"a1"),
   495 => (x"e2",x"ff",x"c3",x"87"),
   496 => (x"c8",x"49",x"bf",x"97"),
   497 => (x"e1",x"ff",x"c3",x"31"),
   498 => (x"a1",x"4a",x"bf",x"97"),
   499 => (x"c7",x"31",x"c5",x"49"),
   500 => (x"29",x"c9",x"81",x"ff"),
   501 => (x"59",x"fc",x"cb",x"c4"),
   502 => (x"97",x"e7",x"ff",x"c3"),
   503 => (x"32",x"c8",x"4a",x"bf"),
   504 => (x"97",x"e6",x"ff",x"c3"),
   505 => (x"4a",x"a2",x"4b",x"bf"),
   506 => (x"6e",x"92",x"66",x"c4"),
   507 => (x"f8",x"cb",x"c4",x"82"),
   508 => (x"f0",x"cb",x"c4",x"5a"),
   509 => (x"c4",x"78",x"c0",x"48"),
   510 => (x"72",x"48",x"ec",x"cb"),
   511 => (x"cb",x"c4",x"78",x"a1"),
   512 => (x"cb",x"c4",x"48",x"fc"),
   513 => (x"c4",x"78",x"bf",x"f0"),
   514 => (x"c4",x"48",x"c0",x"cc"),
   515 => (x"78",x"bf",x"f4",x"cb"),
   516 => (x"bf",x"d8",x"c7",x"c4"),
   517 => (x"87",x"c9",x"c0",x"02"),
   518 => (x"30",x"c4",x"48",x"74"),
   519 => (x"c9",x"c0",x"7e",x"70"),
   520 => (x"f8",x"cb",x"c4",x"87"),
   521 => (x"30",x"c4",x"48",x"bf"),
   522 => (x"c7",x"c4",x"7e",x"70"),
   523 => (x"78",x"6e",x"48",x"dc"),
   524 => (x"8e",x"f8",x"48",x"c1"),
   525 => (x"4c",x"26",x"4d",x"26"),
   526 => (x"4f",x"26",x"4b",x"26"),
   527 => (x"5c",x"5b",x"5e",x"0e"),
   528 => (x"4a",x"71",x"0e",x"5d"),
   529 => (x"bf",x"d8",x"c7",x"c4"),
   530 => (x"72",x"87",x"cb",x"02"),
   531 => (x"72",x"2b",x"c7",x"4b"),
   532 => (x"9d",x"ff",x"c1",x"4d"),
   533 => (x"4b",x"72",x"87",x"c9"),
   534 => (x"4d",x"72",x"2b",x"c8"),
   535 => (x"c4",x"9d",x"ff",x"c3"),
   536 => (x"83",x"bf",x"e8",x"cb"),
   537 => (x"bf",x"c8",x"c2",x"c1"),
   538 => (x"87",x"d9",x"02",x"ab"),
   539 => (x"5b",x"cc",x"c2",x"c1"),
   540 => (x"1e",x"d0",x"ff",x"c3"),
   541 => (x"c5",x"f1",x"49",x"73"),
   542 => (x"70",x"86",x"c4",x"87"),
   543 => (x"87",x"c5",x"05",x"98"),
   544 => (x"e6",x"c0",x"48",x"c0"),
   545 => (x"d8",x"c7",x"c4",x"87"),
   546 => (x"87",x"d2",x"02",x"bf"),
   547 => (x"91",x"c4",x"49",x"75"),
   548 => (x"81",x"d0",x"ff",x"c3"),
   549 => (x"ff",x"cf",x"4c",x"69"),
   550 => (x"9c",x"ff",x"ff",x"ff"),
   551 => (x"49",x"75",x"87",x"cb"),
   552 => (x"ff",x"c3",x"91",x"c2"),
   553 => (x"69",x"9f",x"81",x"d0"),
   554 => (x"26",x"48",x"74",x"4c"),
   555 => (x"26",x"4c",x"26",x"4d"),
   556 => (x"0e",x"4f",x"26",x"4b"),
   557 => (x"5d",x"5c",x"5b",x"5e"),
   558 => (x"cc",x"86",x"f0",x"0e"),
   559 => (x"66",x"c8",x"59",x"a6"),
   560 => (x"c0",x"87",x"c5",x"05"),
   561 => (x"87",x"c4",x"c4",x"48"),
   562 => (x"c8",x"48",x"66",x"c8"),
   563 => (x"48",x"7e",x"70",x"80"),
   564 => (x"e0",x"c0",x"78",x"c0"),
   565 => (x"87",x"c8",x"02",x"66"),
   566 => (x"97",x"66",x"e0",x"c0"),
   567 => (x"87",x"c5",x"05",x"bf"),
   568 => (x"e7",x"c3",x"48",x"c0"),
   569 => (x"c1",x"1e",x"c0",x"87"),
   570 => (x"c2",x"d1",x"49",x"49"),
   571 => (x"70",x"86",x"c4",x"87"),
   572 => (x"c0",x"02",x"9c",x"4c"),
   573 => (x"c7",x"c4",x"87",x"fe"),
   574 => (x"e0",x"c0",x"4a",x"e0"),
   575 => (x"dd",x"ff",x"49",x"66"),
   576 => (x"98",x"70",x"87",x"e7"),
   577 => (x"87",x"ec",x"c0",x"02"),
   578 => (x"e0",x"c0",x"4a",x"74"),
   579 => (x"4b",x"cb",x"49",x"66"),
   580 => (x"87",x"ca",x"de",x"ff"),
   581 => (x"db",x"02",x"98",x"70"),
   582 => (x"74",x"1e",x"c0",x"87"),
   583 => (x"87",x"c4",x"02",x"9c"),
   584 => (x"87",x"c2",x"4d",x"c0"),
   585 => (x"49",x"75",x"4d",x"c1"),
   586 => (x"c4",x"87",x"c4",x"d0"),
   587 => (x"9c",x"4c",x"70",x"86"),
   588 => (x"87",x"c2",x"ff",x"05"),
   589 => (x"c2",x"02",x"9c",x"74"),
   590 => (x"a4",x"dc",x"87",x"d0"),
   591 => (x"69",x"48",x"6e",x"49"),
   592 => (x"49",x"a4",x"da",x"78"),
   593 => (x"c4",x"48",x"66",x"c8"),
   594 => (x"58",x"a6",x"c8",x"80"),
   595 => (x"c4",x"48",x"69",x"9f"),
   596 => (x"c4",x"78",x"08",x"66"),
   597 => (x"02",x"bf",x"d8",x"c7"),
   598 => (x"a4",x"d4",x"87",x"d2"),
   599 => (x"49",x"69",x"9f",x"49"),
   600 => (x"99",x"ff",x"ff",x"c0"),
   601 => (x"30",x"d0",x"48",x"71"),
   602 => (x"87",x"c5",x"58",x"a6"),
   603 => (x"c0",x"48",x"a6",x"cc"),
   604 => (x"48",x"66",x"cc",x"78"),
   605 => (x"80",x"bf",x"66",x"c4"),
   606 => (x"78",x"08",x"66",x"c4"),
   607 => (x"c0",x"48",x"66",x"c8"),
   608 => (x"49",x"66",x"c8",x"78"),
   609 => (x"66",x"c4",x"81",x"cc"),
   610 => (x"66",x"c8",x"79",x"bf"),
   611 => (x"c0",x"81",x"d0",x"49"),
   612 => (x"66",x"c4",x"4d",x"79"),
   613 => (x"4a",x"66",x"c8",x"4c"),
   614 => (x"49",x"75",x"82",x"d4"),
   615 => (x"a1",x"72",x"91",x"c8"),
   616 => (x"6c",x"41",x"c0",x"49"),
   617 => (x"c6",x"85",x"c1",x"79"),
   618 => (x"ff",x"04",x"ad",x"b7"),
   619 => (x"bf",x"6e",x"87",x"e7"),
   620 => (x"72",x"2a",x"c9",x"4a"),
   621 => (x"4a",x"f0",x"c0",x"49"),
   622 => (x"87",x"e3",x"dc",x"ff"),
   623 => (x"66",x"c8",x"4a",x"70"),
   624 => (x"81",x"c4",x"c1",x"49"),
   625 => (x"48",x"c1",x"79",x"72"),
   626 => (x"48",x"c0",x"87",x"c2"),
   627 => (x"4d",x"26",x"8e",x"f0"),
   628 => (x"4b",x"26",x"4c",x"26"),
   629 => (x"5e",x"0e",x"4f",x"26"),
   630 => (x"0e",x"5d",x"5c",x"5b"),
   631 => (x"66",x"d0",x"4c",x"71"),
   632 => (x"02",x"9c",x"74",x"4d"),
   633 => (x"c8",x"87",x"c2",x"c1"),
   634 => (x"02",x"69",x"49",x"a4"),
   635 => (x"6c",x"87",x"fa",x"c0"),
   636 => (x"b9",x"75",x"85",x"49"),
   637 => (x"bf",x"d4",x"c7",x"c4"),
   638 => (x"72",x"ba",x"ff",x"4a"),
   639 => (x"02",x"99",x"71",x"99"),
   640 => (x"c4",x"87",x"e4",x"c0"),
   641 => (x"49",x"6b",x"4b",x"a4"),
   642 => (x"70",x"87",x"f1",x"f8"),
   643 => (x"d0",x"c7",x"c4",x"7b"),
   644 => (x"81",x"6c",x"49",x"bf"),
   645 => (x"b9",x"75",x"7c",x"71"),
   646 => (x"bf",x"d4",x"c7",x"c4"),
   647 => (x"72",x"ba",x"ff",x"4a"),
   648 => (x"05",x"99",x"71",x"99"),
   649 => (x"75",x"87",x"dc",x"ff"),
   650 => (x"26",x"4d",x"26",x"7c"),
   651 => (x"26",x"4b",x"26",x"4c"),
   652 => (x"1e",x"73",x"1e",x"4f"),
   653 => (x"02",x"9b",x"4b",x"71"),
   654 => (x"a3",x"c8",x"87",x"c7"),
   655 => (x"c5",x"05",x"69",x"49"),
   656 => (x"c0",x"48",x"c0",x"87"),
   657 => (x"cb",x"c4",x"87",x"f6"),
   658 => (x"c4",x"49",x"bf",x"ec"),
   659 => (x"4a",x"6a",x"4a",x"a3"),
   660 => (x"c7",x"c4",x"8a",x"c2"),
   661 => (x"72",x"92",x"bf",x"d0"),
   662 => (x"c7",x"c4",x"49",x"a1"),
   663 => (x"6b",x"4a",x"bf",x"d4"),
   664 => (x"49",x"a1",x"72",x"9a"),
   665 => (x"59",x"cc",x"c2",x"c1"),
   666 => (x"71",x"1e",x"66",x"c8"),
   667 => (x"c4",x"87",x"cf",x"e9"),
   668 => (x"05",x"98",x"70",x"86"),
   669 => (x"48",x"c0",x"87",x"c4"),
   670 => (x"48",x"c1",x"87",x"c2"),
   671 => (x"4f",x"26",x"4b",x"26"),
   672 => (x"71",x"1e",x"73",x"1e"),
   673 => (x"c7",x"02",x"9b",x"4b"),
   674 => (x"49",x"a3",x"c8",x"87"),
   675 => (x"87",x"c5",x"05",x"69"),
   676 => (x"f6",x"c0",x"48",x"c0"),
   677 => (x"ec",x"cb",x"c4",x"87"),
   678 => (x"a3",x"c4",x"49",x"bf"),
   679 => (x"c2",x"4a",x"6a",x"4a"),
   680 => (x"d0",x"c7",x"c4",x"8a"),
   681 => (x"a1",x"72",x"92",x"bf"),
   682 => (x"d4",x"c7",x"c4",x"49"),
   683 => (x"9a",x"6b",x"4a",x"bf"),
   684 => (x"c1",x"49",x"a1",x"72"),
   685 => (x"c8",x"59",x"cc",x"c2"),
   686 => (x"e4",x"71",x"1e",x"66"),
   687 => (x"86",x"c4",x"87",x"f1"),
   688 => (x"c4",x"05",x"98",x"70"),
   689 => (x"c2",x"48",x"c0",x"87"),
   690 => (x"26",x"48",x"c1",x"87"),
   691 => (x"0e",x"4f",x"26",x"4b"),
   692 => (x"5d",x"5c",x"5b",x"5e"),
   693 => (x"71",x"86",x"f8",x"0e"),
   694 => (x"48",x"a6",x"c4",x"7e"),
   695 => (x"ff",x"c1",x"78",x"ff"),
   696 => (x"ff",x"ff",x"ff",x"ff"),
   697 => (x"6e",x"4b",x"c0",x"4d"),
   698 => (x"73",x"82",x"d4",x"4a"),
   699 => (x"72",x"91",x"c8",x"49"),
   700 => (x"66",x"d8",x"49",x"a1"),
   701 => (x"c0",x"8c",x"69",x"4c"),
   702 => (x"cb",x"04",x"ac",x"b7"),
   703 => (x"ac",x"b7",x"75",x"87"),
   704 => (x"c8",x"87",x"c5",x"03"),
   705 => (x"4d",x"74",x"5b",x"a6"),
   706 => (x"b7",x"c6",x"83",x"c1"),
   707 => (x"d6",x"ff",x"04",x"ab"),
   708 => (x"48",x"66",x"c4",x"87"),
   709 => (x"4d",x"26",x"8e",x"f8"),
   710 => (x"4b",x"26",x"4c",x"26"),
   711 => (x"5e",x"0e",x"4f",x"26"),
   712 => (x"0e",x"5d",x"5c",x"5b"),
   713 => (x"7e",x"71",x"86",x"f0"),
   714 => (x"c1",x"48",x"a6",x"c4"),
   715 => (x"ff",x"ff",x"ff",x"ff"),
   716 => (x"80",x"c4",x"78",x"ff"),
   717 => (x"4d",x"c0",x"78",x"ff"),
   718 => (x"4b",x"6e",x"4c",x"c0"),
   719 => (x"4a",x"74",x"83",x"d4"),
   720 => (x"a2",x"73",x"92",x"c8"),
   721 => (x"c8",x"49",x"75",x"4a"),
   722 => (x"49",x"a1",x"73",x"91"),
   723 => (x"88",x"69",x"48",x"6a"),
   724 => (x"a6",x"d0",x"49",x"70"),
   725 => (x"02",x"ad",x"74",x"59"),
   726 => (x"66",x"cc",x"87",x"d2"),
   727 => (x"a8",x"66",x"c4",x"48"),
   728 => (x"cc",x"87",x"c9",x"03"),
   729 => (x"a6",x"c4",x"5c",x"a6"),
   730 => (x"78",x"66",x"cc",x"48"),
   731 => (x"b7",x"c6",x"84",x"c1"),
   732 => (x"c5",x"ff",x"04",x"ac"),
   733 => (x"c6",x"85",x"c1",x"87"),
   734 => (x"fe",x"04",x"ad",x"b7"),
   735 => (x"66",x"c8",x"87",x"fa"),
   736 => (x"26",x"8e",x"f0",x"48"),
   737 => (x"26",x"4c",x"26",x"4d"),
   738 => (x"0e",x"4f",x"26",x"4b"),
   739 => (x"5d",x"5c",x"5b",x"5e"),
   740 => (x"71",x"86",x"ec",x"0e"),
   741 => (x"66",x"e4",x"c0",x"4b"),
   742 => (x"c8",x"28",x"c9",x"48"),
   743 => (x"c7",x"c4",x"58",x"a6"),
   744 => (x"ff",x"4a",x"bf",x"d4"),
   745 => (x"c4",x"48",x"72",x"ba"),
   746 => (x"a6",x"cc",x"98",x"66"),
   747 => (x"02",x"9b",x"73",x"58"),
   748 => (x"c8",x"87",x"c1",x"c3"),
   749 => (x"02",x"69",x"49",x"a3"),
   750 => (x"72",x"87",x"f9",x"c2"),
   751 => (x"d4",x"98",x"6b",x"48"),
   752 => (x"a3",x"c4",x"58",x"a6"),
   753 => (x"c8",x"7e",x"6c",x"4c"),
   754 => (x"66",x"d0",x"48",x"66"),
   755 => (x"87",x"c6",x"05",x"a8"),
   756 => (x"c2",x"7b",x"66",x"c4"),
   757 => (x"66",x"c8",x"87",x"cc"),
   758 => (x"fb",x"49",x"73",x"1e"),
   759 => (x"86",x"c4",x"87",x"f1"),
   760 => (x"b7",x"c0",x"4d",x"70"),
   761 => (x"87",x"d0",x"04",x"ad"),
   762 => (x"75",x"4a",x"a3",x"d4"),
   763 => (x"72",x"91",x"c8",x"49"),
   764 => (x"7b",x"21",x"49",x"a1"),
   765 => (x"87",x"c7",x"7c",x"69"),
   766 => (x"a3",x"cc",x"7b",x"c0"),
   767 => (x"c4",x"7c",x"69",x"49"),
   768 => (x"88",x"6b",x"48",x"66"),
   769 => (x"d0",x"58",x"a6",x"c8"),
   770 => (x"49",x"73",x"1e",x"66"),
   771 => (x"c4",x"87",x"c0",x"fb"),
   772 => (x"c1",x"4d",x"70",x"86"),
   773 => (x"c8",x"49",x"a3",x"c4"),
   774 => (x"78",x"69",x"48",x"a6"),
   775 => (x"c8",x"48",x"66",x"d0"),
   776 => (x"c0",x"06",x"a8",x"66"),
   777 => (x"b7",x"c0",x"87",x"f2"),
   778 => (x"eb",x"c0",x"04",x"ad"),
   779 => (x"48",x"a6",x"cc",x"87"),
   780 => (x"75",x"78",x"a3",x"d4"),
   781 => (x"cc",x"91",x"c8",x"49"),
   782 => (x"66",x"d0",x"81",x"66"),
   783 => (x"70",x"88",x"69",x"48"),
   784 => (x"a9",x"66",x"c8",x"49"),
   785 => (x"73",x"87",x"d1",x"06"),
   786 => (x"87",x"d2",x"fb",x"49"),
   787 => (x"91",x"c8",x"49",x"70"),
   788 => (x"d0",x"81",x"66",x"cc"),
   789 => (x"79",x"6e",x"41",x"66"),
   790 => (x"73",x"1e",x"66",x"c4"),
   791 => (x"87",x"f6",x"f5",x"49"),
   792 => (x"ff",x"c3",x"86",x"c4"),
   793 => (x"49",x"73",x"1e",x"d0"),
   794 => (x"c4",x"87",x"c6",x"f7"),
   795 => (x"49",x"a3",x"d0",x"86"),
   796 => (x"79",x"66",x"e4",x"c0"),
   797 => (x"4d",x"26",x"8e",x"ec"),
   798 => (x"4b",x"26",x"4c",x"26"),
   799 => (x"73",x"1e",x"4f",x"26"),
   800 => (x"9b",x"4b",x"71",x"1e"),
   801 => (x"87",x"e4",x"c0",x"02"),
   802 => (x"5b",x"c0",x"cc",x"c4"),
   803 => (x"8a",x"c2",x"4a",x"73"),
   804 => (x"bf",x"d0",x"c7",x"c4"),
   805 => (x"cb",x"c4",x"92",x"49"),
   806 => (x"72",x"48",x"bf",x"ec"),
   807 => (x"c4",x"cc",x"c4",x"80"),
   808 => (x"c4",x"48",x"71",x"58"),
   809 => (x"e0",x"c7",x"c4",x"30"),
   810 => (x"87",x"ed",x"c0",x"58"),
   811 => (x"48",x"fc",x"cb",x"c4"),
   812 => (x"bf",x"f0",x"cb",x"c4"),
   813 => (x"c0",x"cc",x"c4",x"78"),
   814 => (x"f4",x"cb",x"c4",x"48"),
   815 => (x"c7",x"c4",x"78",x"bf"),
   816 => (x"c9",x"02",x"bf",x"d8"),
   817 => (x"d0",x"c7",x"c4",x"87"),
   818 => (x"31",x"c4",x"49",x"bf"),
   819 => (x"cb",x"c4",x"87",x"c7"),
   820 => (x"c4",x"49",x"bf",x"f8"),
   821 => (x"e0",x"c7",x"c4",x"31"),
   822 => (x"26",x"4b",x"26",x"59"),
   823 => (x"cb",x"c4",x"1e",x"4f"),
   824 => (x"c4",x"49",x"bf",x"fc"),
   825 => (x"a9",x"bf",x"f0",x"cb"),
   826 => (x"c0",x"87",x"c4",x"05"),
   827 => (x"71",x"87",x"c2",x"4a"),
   828 => (x"26",x"48",x"72",x"4a"),
   829 => (x"5b",x"5e",x"0e",x"4f"),
   830 => (x"4a",x"71",x"0e",x"5c"),
   831 => (x"9a",x"72",x"4b",x"c0"),
   832 => (x"87",x"e0",x"c0",x"02"),
   833 => (x"9f",x"49",x"a2",x"da"),
   834 => (x"c7",x"c4",x"4b",x"69"),
   835 => (x"cf",x"02",x"bf",x"d8"),
   836 => (x"49",x"a2",x"d4",x"87"),
   837 => (x"4c",x"49",x"69",x"9f"),
   838 => (x"9c",x"ff",x"ff",x"c0"),
   839 => (x"87",x"c2",x"34",x"d0"),
   840 => (x"b3",x"74",x"4c",x"c0"),
   841 => (x"d5",x"fd",x"49",x"73"),
   842 => (x"26",x"4c",x"26",x"87"),
   843 => (x"0e",x"4f",x"26",x"4b"),
   844 => (x"5d",x"5c",x"5b",x"5e"),
   845 => (x"c8",x"86",x"f0",x"0e"),
   846 => (x"ff",x"cf",x"59",x"a6"),
   847 => (x"4c",x"f8",x"ff",x"ff"),
   848 => (x"66",x"c4",x"7e",x"c0"),
   849 => (x"c3",x"87",x"d8",x"02"),
   850 => (x"c0",x"48",x"cc",x"ff"),
   851 => (x"c4",x"ff",x"c3",x"78"),
   852 => (x"c0",x"cc",x"c4",x"48"),
   853 => (x"ff",x"c3",x"78",x"bf"),
   854 => (x"cb",x"c4",x"48",x"c8"),
   855 => (x"c4",x"78",x"bf",x"fc"),
   856 => (x"c0",x"48",x"ed",x"c7"),
   857 => (x"dc",x"c7",x"c4",x"50"),
   858 => (x"ff",x"c3",x"49",x"bf"),
   859 => (x"71",x"4a",x"bf",x"cc"),
   860 => (x"cc",x"c4",x"03",x"aa"),
   861 => (x"cf",x"49",x"72",x"87"),
   862 => (x"ea",x"c0",x"05",x"99"),
   863 => (x"c8",x"c2",x"c1",x"87"),
   864 => (x"c4",x"ff",x"c3",x"48"),
   865 => (x"ff",x"c3",x"78",x"bf"),
   866 => (x"ff",x"c3",x"1e",x"d0"),
   867 => (x"c3",x"49",x"bf",x"c4"),
   868 => (x"c1",x"48",x"c4",x"ff"),
   869 => (x"ff",x"71",x"78",x"a1"),
   870 => (x"c4",x"87",x"e3",x"dc"),
   871 => (x"e4",x"fc",x"c0",x"86"),
   872 => (x"d0",x"ff",x"c3",x"48"),
   873 => (x"c0",x"87",x"cc",x"78"),
   874 => (x"48",x"bf",x"e4",x"fc"),
   875 => (x"c0",x"80",x"e0",x"c0"),
   876 => (x"c3",x"58",x"e8",x"fc"),
   877 => (x"48",x"bf",x"cc",x"ff"),
   878 => (x"ff",x"c3",x"80",x"c1"),
   879 => (x"24",x"27",x"58",x"d0"),
   880 => (x"bf",x"00",x"00",x"0f"),
   881 => (x"9d",x"4d",x"bf",x"97"),
   882 => (x"87",x"e5",x"c2",x"02"),
   883 => (x"02",x"ad",x"e5",x"c3"),
   884 => (x"c0",x"87",x"de",x"c2"),
   885 => (x"4b",x"bf",x"e4",x"fc"),
   886 => (x"11",x"49",x"a3",x"cb"),
   887 => (x"05",x"ac",x"cf",x"4c"),
   888 => (x"75",x"87",x"d2",x"c1"),
   889 => (x"c1",x"99",x"df",x"49"),
   890 => (x"c4",x"91",x"cd",x"89"),
   891 => (x"c1",x"81",x"e0",x"c7"),
   892 => (x"51",x"12",x"4a",x"a3"),
   893 => (x"12",x"4a",x"a3",x"c3"),
   894 => (x"4a",x"a3",x"c5",x"51"),
   895 => (x"a3",x"c7",x"51",x"12"),
   896 => (x"c9",x"51",x"12",x"4a"),
   897 => (x"51",x"12",x"4a",x"a3"),
   898 => (x"12",x"4a",x"a3",x"ce"),
   899 => (x"4a",x"a3",x"d0",x"51"),
   900 => (x"a3",x"d2",x"51",x"12"),
   901 => (x"d4",x"51",x"12",x"4a"),
   902 => (x"51",x"12",x"4a",x"a3"),
   903 => (x"12",x"4a",x"a3",x"d6"),
   904 => (x"4a",x"a3",x"d8",x"51"),
   905 => (x"a3",x"dc",x"51",x"12"),
   906 => (x"de",x"51",x"12",x"4a"),
   907 => (x"51",x"12",x"4a",x"a3"),
   908 => (x"fc",x"c0",x"7e",x"c1"),
   909 => (x"c8",x"49",x"74",x"87"),
   910 => (x"ed",x"c0",x"05",x"99"),
   911 => (x"d0",x"49",x"74",x"87"),
   912 => (x"87",x"d3",x"05",x"99"),
   913 => (x"02",x"66",x"e0",x"c0"),
   914 => (x"73",x"87",x"cc",x"c0"),
   915 => (x"66",x"e0",x"c0",x"49"),
   916 => (x"02",x"98",x"70",x"0f"),
   917 => (x"6e",x"87",x"d3",x"c0"),
   918 => (x"87",x"c6",x"c0",x"05"),
   919 => (x"48",x"e0",x"c7",x"c4"),
   920 => (x"fc",x"c0",x"50",x"c0"),
   921 => (x"c2",x"48",x"bf",x"e4"),
   922 => (x"c7",x"c4",x"87",x"e9"),
   923 => (x"50",x"c0",x"48",x"ed"),
   924 => (x"dc",x"c7",x"c4",x"7e"),
   925 => (x"ff",x"c3",x"49",x"bf"),
   926 => (x"71",x"4a",x"bf",x"cc"),
   927 => (x"f4",x"fb",x"04",x"aa"),
   928 => (x"ff",x"ff",x"cf",x"87"),
   929 => (x"c4",x"4c",x"f8",x"ff"),
   930 => (x"05",x"bf",x"c0",x"cc"),
   931 => (x"c4",x"87",x"c8",x"c0"),
   932 => (x"02",x"bf",x"d8",x"c7"),
   933 => (x"c3",x"87",x"fa",x"c1"),
   934 => (x"49",x"bf",x"c8",x"ff"),
   935 => (x"c3",x"87",x"dd",x"e6"),
   936 => (x"c4",x"58",x"cc",x"ff"),
   937 => (x"ff",x"c3",x"48",x"a6"),
   938 => (x"c4",x"78",x"bf",x"c8"),
   939 => (x"02",x"bf",x"d8",x"c7"),
   940 => (x"c4",x"87",x"db",x"c0"),
   941 => (x"99",x"74",x"49",x"66"),
   942 => (x"c0",x"02",x"a9",x"74"),
   943 => (x"a6",x"c8",x"87",x"c8"),
   944 => (x"c0",x"78",x"c0",x"48"),
   945 => (x"a6",x"c8",x"87",x"e7"),
   946 => (x"c0",x"78",x"c1",x"48"),
   947 => (x"66",x"c4",x"87",x"df"),
   948 => (x"f8",x"ff",x"cf",x"49"),
   949 => (x"c0",x"02",x"a9",x"99"),
   950 => (x"a6",x"cc",x"87",x"c8"),
   951 => (x"c0",x"78",x"c0",x"48"),
   952 => (x"a6",x"cc",x"87",x"c5"),
   953 => (x"c8",x"78",x"c1",x"48"),
   954 => (x"66",x"cc",x"48",x"a6"),
   955 => (x"05",x"66",x"c8",x"78"),
   956 => (x"c4",x"87",x"de",x"c0"),
   957 => (x"89",x"c2",x"49",x"66"),
   958 => (x"bf",x"d0",x"c7",x"c4"),
   959 => (x"ec",x"cb",x"c4",x"91"),
   960 => (x"80",x"71",x"48",x"bf"),
   961 => (x"58",x"c8",x"ff",x"c3"),
   962 => (x"48",x"cc",x"ff",x"c3"),
   963 => (x"d4",x"f9",x"78",x"c0"),
   964 => (x"cf",x"48",x"c0",x"87"),
   965 => (x"f8",x"ff",x"ff",x"ff"),
   966 => (x"26",x"8e",x"f0",x"4c"),
   967 => (x"26",x"4c",x"26",x"4d"),
   968 => (x"00",x"4f",x"26",x"4b"),
   969 => (x"00",x"00",x"00",x"00"),
   970 => (x"5c",x"5b",x"5e",x"0e"),
   971 => (x"86",x"fc",x"0e",x"5d"),
   972 => (x"49",x"6e",x"7e",x"71"),
   973 => (x"c0",x"87",x"c7",x"f5"),
   974 => (x"49",x"49",x"c1",x"1e"),
   975 => (x"c4",x"87",x"f0",x"f7"),
   976 => (x"9a",x"4a",x"70",x"86"),
   977 => (x"87",x"c6",x"c1",x"02"),
   978 => (x"9f",x"49",x"a2",x"da"),
   979 => (x"c7",x"c4",x"4b",x"69"),
   980 => (x"cf",x"02",x"bf",x"d8"),
   981 => (x"49",x"a2",x"d4",x"87"),
   982 => (x"4c",x"49",x"69",x"9f"),
   983 => (x"9c",x"ff",x"ff",x"c0"),
   984 => (x"87",x"c2",x"34",x"d0"),
   985 => (x"a3",x"74",x"4c",x"c0"),
   986 => (x"ab",x"66",x"d4",x"4b"),
   987 => (x"c1",x"87",x"c4",x"05"),
   988 => (x"c0",x"87",x"dd",x"48"),
   989 => (x"02",x"9a",x"72",x"1e"),
   990 => (x"4d",x"c0",x"87",x"c4"),
   991 => (x"4d",x"c1",x"87",x"c2"),
   992 => (x"ea",x"f6",x"49",x"75"),
   993 => (x"70",x"86",x"c4",x"87"),
   994 => (x"fe",x"05",x"9a",x"4a"),
   995 => (x"48",x"c0",x"87",x"fa"),
   996 => (x"4d",x"26",x"8e",x"fc"),
   997 => (x"4b",x"26",x"4c",x"26"),
   998 => (x"5e",x"0e",x"4f",x"26"),
   999 => (x"0e",x"5d",x"5c",x"5b"),
  1000 => (x"a6",x"c8",x"86",x"f4"),
  1001 => (x"02",x"66",x"c4",x"59"),
  1002 => (x"c4",x"48",x"87",x"c9"),
  1003 => (x"a8",x"bf",x"f0",x"cb"),
  1004 => (x"c1",x"87",x"c5",x"05"),
  1005 => (x"87",x"f7",x"c2",x"48"),
  1006 => (x"c2",x"49",x"66",x"c4"),
  1007 => (x"d0",x"c7",x"c4",x"89"),
  1008 => (x"cb",x"c4",x"91",x"bf"),
  1009 => (x"c3",x"81",x"bf",x"ec"),
  1010 => (x"71",x"1e",x"d0",x"ff"),
  1011 => (x"87",x"ee",x"d3",x"ff"),
  1012 => (x"98",x"70",x"86",x"c4"),
  1013 => (x"c0",x"87",x"c5",x"05"),
  1014 => (x"87",x"d3",x"c2",x"48"),
  1015 => (x"4c",x"d0",x"ff",x"c3"),
  1016 => (x"6c",x"97",x"7e",x"c0"),
  1017 => (x"58",x"a6",x"cc",x"48"),
  1018 => (x"c1",x"02",x"98",x"70"),
  1019 => (x"c3",x"48",x"87",x"ef"),
  1020 => (x"c1",x"02",x"a8",x"e5"),
  1021 => (x"a4",x"cb",x"87",x"e7"),
  1022 => (x"49",x"69",x"97",x"49"),
  1023 => (x"c1",x"02",x"99",x"d0"),
  1024 => (x"4a",x"74",x"87",x"db"),
  1025 => (x"49",x"fc",x"c1",x"c1"),
  1026 => (x"c1",x"ff",x"4b",x"c8"),
  1027 => (x"98",x"70",x"87",x"f6"),
  1028 => (x"87",x"c9",x"c1",x"05"),
  1029 => (x"c4",x"7e",x"a4",x"da"),
  1030 => (x"02",x"bf",x"d8",x"c7"),
  1031 => (x"a4",x"d4",x"87",x"cf"),
  1032 => (x"49",x"69",x"9f",x"49"),
  1033 => (x"ff",x"ff",x"c0",x"4d"),
  1034 => (x"c2",x"35",x"d0",x"9d"),
  1035 => (x"6e",x"4d",x"c0",x"87"),
  1036 => (x"75",x"49",x"bf",x"9f"),
  1037 => (x"59",x"a6",x"cc",x"81"),
  1038 => (x"fd",x"49",x"66",x"c8"),
  1039 => (x"98",x"70",x"87",x"dc"),
  1040 => (x"c4",x"87",x"d4",x"02"),
  1041 => (x"66",x"cc",x"1e",x"66"),
  1042 => (x"87",x"dc",x"fb",x"49"),
  1043 => (x"98",x"70",x"86",x"c4"),
  1044 => (x"c1",x"87",x"c4",x"02"),
  1045 => (x"c0",x"87",x"c2",x"7e"),
  1046 => (x"d2",x"48",x"6e",x"7e"),
  1047 => (x"84",x"e0",x"c0",x"87"),
  1048 => (x"80",x"c1",x"48",x"6e"),
  1049 => (x"d0",x"48",x"7e",x"70"),
  1050 => (x"f5",x"fd",x"04",x"a8"),
  1051 => (x"f4",x"48",x"c0",x"87"),
  1052 => (x"26",x"4d",x"26",x"8e"),
  1053 => (x"26",x"4b",x"26",x"4c"),
  1054 => (x"00",x"00",x"00",x"4f"),
  1055 => (x"20",x"20",x"2e",x"2e"),
  1056 => (x"20",x"20",x"20",x"20"),
  1057 => (x"00",x"20",x"20",x"20"),
  1058 => (x"ff",x"ff",x"ff",x"ff"),
  1059 => (x"00",x"00",x"10",x"94"),
  1060 => (x"00",x"00",x"10",x"a0"),
  1061 => (x"33",x"54",x"41",x"46"),
  1062 => (x"20",x"20",x"20",x"32"),
  1063 => (x"00",x"00",x"00",x"00"),
  1064 => (x"31",x"54",x"41",x"46"),
  1065 => (x"20",x"20",x"20",x"36"),
  1066 => (x"d0",x"ff",x"1e",x"00"),
  1067 => (x"78",x"e0",x"c0",x"48"),
  1068 => (x"c2",x"1e",x"4f",x"26"),
  1069 => (x"70",x"87",x"d9",x"d2"),
  1070 => (x"c6",x"02",x"99",x"49"),
  1071 => (x"a9",x"fb",x"c0",x"87"),
  1072 => (x"71",x"87",x"f0",x"05"),
  1073 => (x"0e",x"4f",x"26",x"48"),
  1074 => (x"0e",x"5c",x"5b",x"5e"),
  1075 => (x"4c",x"c0",x"4b",x"71"),
  1076 => (x"87",x"fc",x"d1",x"c2"),
  1077 => (x"02",x"99",x"49",x"70"),
  1078 => (x"c0",x"87",x"fa",x"c0"),
  1079 => (x"c0",x"02",x"a9",x"ec"),
  1080 => (x"fb",x"c0",x"87",x"f3"),
  1081 => (x"ec",x"c0",x"02",x"a9"),
  1082 => (x"b7",x"66",x"cc",x"87"),
  1083 => (x"87",x"c7",x"03",x"ac"),
  1084 => (x"c2",x"02",x"66",x"d0"),
  1085 => (x"71",x"53",x"71",x"87"),
  1086 => (x"87",x"c2",x"02",x"99"),
  1087 => (x"d1",x"c2",x"84",x"c1"),
  1088 => (x"49",x"70",x"87",x"ce"),
  1089 => (x"87",x"cd",x"02",x"99"),
  1090 => (x"02",x"a9",x"ec",x"c0"),
  1091 => (x"fb",x"c0",x"87",x"c7"),
  1092 => (x"d4",x"ff",x"05",x"a9"),
  1093 => (x"02",x"66",x"d0",x"87"),
  1094 => (x"97",x"c0",x"87",x"c3"),
  1095 => (x"a9",x"ec",x"c0",x"7b"),
  1096 => (x"74",x"87",x"c4",x"05"),
  1097 => (x"74",x"87",x"c5",x"4a"),
  1098 => (x"8a",x"0a",x"c0",x"4a"),
  1099 => (x"4c",x"26",x"48",x"72"),
  1100 => (x"4f",x"26",x"4b",x"26"),
  1101 => (x"d7",x"d0",x"c2",x"1e"),
  1102 => (x"4a",x"49",x"70",x"87"),
  1103 => (x"04",x"aa",x"f0",x"c0"),
  1104 => (x"f9",x"c0",x"87",x"c9"),
  1105 => (x"87",x"c3",x"01",x"aa"),
  1106 => (x"c1",x"8a",x"f0",x"c0"),
  1107 => (x"c9",x"04",x"aa",x"c1"),
  1108 => (x"aa",x"da",x"c1",x"87"),
  1109 => (x"c0",x"87",x"c3",x"01"),
  1110 => (x"48",x"72",x"8a",x"f7"),
  1111 => (x"5e",x"0e",x"4f",x"26"),
  1112 => (x"0e",x"5d",x"5c",x"5b"),
  1113 => (x"4c",x"71",x"86",x"f8"),
  1114 => (x"d0",x"c2",x"7e",x"c0"),
  1115 => (x"4b",x"c0",x"87",x"c5"),
  1116 => (x"97",x"c4",x"c8",x"c1"),
  1117 => (x"a9",x"c0",x"49",x"bf"),
  1118 => (x"fc",x"87",x"cf",x"04"),
  1119 => (x"83",x"c1",x"87",x"f4"),
  1120 => (x"97",x"c4",x"c8",x"c1"),
  1121 => (x"06",x"ab",x"49",x"bf"),
  1122 => (x"c8",x"c1",x"87",x"f1"),
  1123 => (x"02",x"bf",x"97",x"c4"),
  1124 => (x"ce",x"c2",x"87",x"d0"),
  1125 => (x"49",x"70",x"87",x"fa"),
  1126 => (x"87",x"c6",x"02",x"99"),
  1127 => (x"05",x"a9",x"ec",x"c0"),
  1128 => (x"4b",x"c0",x"87",x"f0"),
  1129 => (x"87",x"e8",x"ce",x"c2"),
  1130 => (x"ce",x"c2",x"4d",x"70"),
  1131 => (x"a6",x"c8",x"87",x"e2"),
  1132 => (x"db",x"ce",x"c2",x"58"),
  1133 => (x"c1",x"4a",x"70",x"87"),
  1134 => (x"49",x"a4",x"c8",x"83"),
  1135 => (x"ad",x"49",x"69",x"97"),
  1136 => (x"c9",x"87",x"da",x"05"),
  1137 => (x"69",x"97",x"49",x"a4"),
  1138 => (x"a9",x"66",x"c4",x"49"),
  1139 => (x"ca",x"87",x"ce",x"05"),
  1140 => (x"69",x"97",x"49",x"a4"),
  1141 => (x"c4",x"05",x"aa",x"49"),
  1142 => (x"d0",x"7e",x"c1",x"87"),
  1143 => (x"ad",x"ec",x"c0",x"87"),
  1144 => (x"c0",x"87",x"c6",x"02"),
  1145 => (x"c4",x"05",x"ad",x"fb"),
  1146 => (x"c1",x"4b",x"c0",x"87"),
  1147 => (x"fe",x"02",x"6e",x"7e"),
  1148 => (x"f4",x"fa",x"87",x"f2"),
  1149 => (x"f8",x"48",x"73",x"87"),
  1150 => (x"26",x"4d",x"26",x"8e"),
  1151 => (x"26",x"4b",x"26",x"4c"),
  1152 => (x"00",x"00",x"00",x"4f"),
  1153 => (x"5b",x"5e",x"0e",x"00"),
  1154 => (x"f4",x"0e",x"5d",x"5c"),
  1155 => (x"ff",x"7e",x"71",x"86"),
  1156 => (x"1e",x"6e",x"4b",x"d4"),
  1157 => (x"49",x"cc",x"cc",x"c4"),
  1158 => (x"87",x"d7",x"da",x"ff"),
  1159 => (x"98",x"70",x"86",x"c4"),
  1160 => (x"87",x"f7",x"c4",x"02"),
  1161 => (x"c1",x"48",x"a6",x"c4"),
  1162 => (x"78",x"bf",x"e8",x"f3"),
  1163 => (x"ed",x"fc",x"49",x"6e"),
  1164 => (x"58",x"a6",x"cc",x"87"),
  1165 => (x"c5",x"05",x"98",x"70"),
  1166 => (x"48",x"a6",x"c8",x"87"),
  1167 => (x"d0",x"ff",x"78",x"c1"),
  1168 => (x"c1",x"78",x"c5",x"48"),
  1169 => (x"66",x"c8",x"7b",x"d5"),
  1170 => (x"c6",x"89",x"c1",x"49"),
  1171 => (x"e0",x"f3",x"c1",x"31"),
  1172 => (x"48",x"4a",x"bf",x"97"),
  1173 => (x"7b",x"70",x"b0",x"71"),
  1174 => (x"c4",x"48",x"d0",x"ff"),
  1175 => (x"c4",x"cc",x"c4",x"78"),
  1176 => (x"d0",x"49",x"bf",x"97"),
  1177 => (x"87",x"d7",x"02",x"99"),
  1178 => (x"d6",x"c1",x"78",x"c5"),
  1179 => (x"c3",x"4a",x"c0",x"7b"),
  1180 => (x"82",x"c1",x"7b",x"ff"),
  1181 => (x"04",x"aa",x"e0",x"c0"),
  1182 => (x"d0",x"ff",x"87",x"f5"),
  1183 => (x"c3",x"78",x"c4",x"48"),
  1184 => (x"d0",x"ff",x"7b",x"ff"),
  1185 => (x"c1",x"78",x"c5",x"48"),
  1186 => (x"7b",x"c1",x"7b",x"d3"),
  1187 => (x"7e",x"73",x"78",x"c4"),
  1188 => (x"c0",x"48",x"66",x"c4"),
  1189 => (x"c2",x"06",x"a8",x"b7"),
  1190 => (x"cc",x"c4",x"87",x"ee"),
  1191 => (x"c4",x"4c",x"bf",x"d4"),
  1192 => (x"88",x"74",x"48",x"66"),
  1193 => (x"74",x"58",x"a6",x"c8"),
  1194 => (x"f7",x"c1",x"02",x"9c"),
  1195 => (x"d0",x"ff",x"c3",x"87"),
  1196 => (x"4b",x"c0",x"c8",x"4d"),
  1197 => (x"ac",x"b7",x"c0",x"8c"),
  1198 => (x"c8",x"87",x"c6",x"03"),
  1199 => (x"c0",x"4b",x"a4",x"c0"),
  1200 => (x"c4",x"cc",x"c4",x"4c"),
  1201 => (x"d0",x"49",x"bf",x"97"),
  1202 => (x"87",x"d1",x"02",x"99"),
  1203 => (x"cc",x"c4",x"1e",x"c0"),
  1204 => (x"dd",x"ff",x"49",x"cc"),
  1205 => (x"86",x"c4",x"87",x"db"),
  1206 => (x"eb",x"c0",x"4a",x"70"),
  1207 => (x"d0",x"ff",x"c3",x"87"),
  1208 => (x"cc",x"cc",x"c4",x"1e"),
  1209 => (x"c8",x"dd",x"ff",x"49"),
  1210 => (x"70",x"86",x"c4",x"87"),
  1211 => (x"48",x"d0",x"ff",x"4a"),
  1212 => (x"6e",x"78",x"c5",x"c8"),
  1213 => (x"78",x"d4",x"c1",x"48"),
  1214 => (x"08",x"6e",x"48",x"15"),
  1215 => (x"05",x"8b",x"c1",x"78"),
  1216 => (x"ff",x"87",x"f5",x"ff"),
  1217 => (x"78",x"c4",x"48",x"d0"),
  1218 => (x"c5",x"05",x"9a",x"72"),
  1219 => (x"c1",x"48",x"c0",x"87"),
  1220 => (x"1e",x"c1",x"87",x"cb"),
  1221 => (x"49",x"cc",x"cc",x"c4"),
  1222 => (x"87",x"fa",x"da",x"ff"),
  1223 => (x"9c",x"74",x"86",x"c4"),
  1224 => (x"87",x"c9",x"fe",x"05"),
  1225 => (x"c0",x"48",x"66",x"c4"),
  1226 => (x"d1",x"06",x"a8",x"b7"),
  1227 => (x"cc",x"cc",x"c4",x"87"),
  1228 => (x"d0",x"78",x"c0",x"48"),
  1229 => (x"f4",x"78",x"c0",x"80"),
  1230 => (x"d8",x"cc",x"c4",x"80"),
  1231 => (x"66",x"c4",x"78",x"bf"),
  1232 => (x"a8",x"b7",x"c0",x"48"),
  1233 => (x"87",x"d2",x"fd",x"01"),
  1234 => (x"d0",x"ff",x"4b",x"6e"),
  1235 => (x"c1",x"78",x"c5",x"48"),
  1236 => (x"7b",x"c0",x"7b",x"d3"),
  1237 => (x"48",x"c1",x"78",x"c4"),
  1238 => (x"c0",x"87",x"c2",x"c0"),
  1239 => (x"26",x"8e",x"f4",x"48"),
  1240 => (x"26",x"4c",x"26",x"4d"),
  1241 => (x"0e",x"4f",x"26",x"4b"),
  1242 => (x"5d",x"5c",x"5b",x"5e"),
  1243 => (x"71",x"86",x"fc",x"0e"),
  1244 => (x"4c",x"4b",x"c0",x"4d"),
  1245 => (x"e8",x"c0",x"04",x"ad"),
  1246 => (x"de",x"c5",x"c1",x"87"),
  1247 => (x"02",x"9c",x"74",x"1e"),
  1248 => (x"4a",x"c0",x"87",x"c4"),
  1249 => (x"4a",x"c1",x"87",x"c2"),
  1250 => (x"e2",x"e6",x"49",x"72"),
  1251 => (x"70",x"86",x"c4",x"87"),
  1252 => (x"6e",x"83",x"c1",x"7e"),
  1253 => (x"75",x"87",x"c2",x"05"),
  1254 => (x"75",x"84",x"c1",x"4b"),
  1255 => (x"d8",x"ff",x"06",x"ab"),
  1256 => (x"fc",x"48",x"6e",x"87"),
  1257 => (x"26",x"4d",x"26",x"8e"),
  1258 => (x"26",x"4b",x"26",x"4c"),
  1259 => (x"5b",x"5e",x"0e",x"4f"),
  1260 => (x"fc",x"0e",x"5d",x"5c"),
  1261 => (x"49",x"4c",x"71",x"86"),
  1262 => (x"cd",x"c4",x"91",x"de"),
  1263 => (x"85",x"71",x"4d",x"e8"),
  1264 => (x"c1",x"02",x"6d",x"97"),
  1265 => (x"cd",x"c4",x"87",x"dd"),
  1266 => (x"74",x"49",x"bf",x"d4"),
  1267 => (x"d6",x"fe",x"71",x"81"),
  1268 => (x"48",x"7e",x"70",x"87"),
  1269 => (x"f3",x"c0",x"02",x"98"),
  1270 => (x"dc",x"cd",x"c4",x"87"),
  1271 => (x"cb",x"4a",x"70",x"4b"),
  1272 => (x"dd",x"f3",x"fe",x"49"),
  1273 => (x"cc",x"4b",x"74",x"87"),
  1274 => (x"fc",x"f3",x"c1",x"93"),
  1275 => (x"c1",x"83",x"c4",x"83"),
  1276 => (x"74",x"7b",x"f0",x"d0"),
  1277 => (x"df",x"c6",x"c1",x"49"),
  1278 => (x"c1",x"7b",x"75",x"87"),
  1279 => (x"bf",x"97",x"e4",x"f3"),
  1280 => (x"cd",x"c4",x"1e",x"49"),
  1281 => (x"d5",x"c2",x"49",x"dc"),
  1282 => (x"86",x"c4",x"87",x"ce"),
  1283 => (x"c6",x"c1",x"49",x"74"),
  1284 => (x"49",x"c0",x"87",x"c6"),
  1285 => (x"87",x"e1",x"c7",x"c1"),
  1286 => (x"48",x"c8",x"cc",x"c4"),
  1287 => (x"49",x"c1",x"78",x"c0"),
  1288 => (x"fc",x"87",x"c4",x"de"),
  1289 => (x"26",x"4d",x"26",x"8e"),
  1290 => (x"26",x"4b",x"26",x"4c"),
  1291 => (x"00",x"00",x"00",x"4f"),
  1292 => (x"64",x"61",x"6f",x"4c"),
  1293 => (x"2e",x"67",x"6e",x"69"),
  1294 => (x"1e",x"00",x"2e",x"2e"),
  1295 => (x"4a",x"71",x"1e",x"73"),
  1296 => (x"d4",x"cd",x"c4",x"49"),
  1297 => (x"fc",x"71",x"81",x"bf"),
  1298 => (x"4b",x"70",x"87",x"dd"),
  1299 => (x"87",x"c4",x"02",x"9b"),
  1300 => (x"87",x"e1",x"e2",x"49"),
  1301 => (x"48",x"d4",x"cd",x"c4"),
  1302 => (x"49",x"c1",x"78",x"c0"),
  1303 => (x"26",x"87",x"c8",x"dd"),
  1304 => (x"1e",x"4f",x"26",x"4b"),
  1305 => (x"c6",x"c1",x"49",x"c0"),
  1306 => (x"4f",x"26",x"87",x"cf"),
  1307 => (x"49",x"4a",x"71",x"1e"),
  1308 => (x"f3",x"c1",x"91",x"cc"),
  1309 => (x"81",x"c8",x"81",x"fc"),
  1310 => (x"cc",x"c4",x"48",x"11"),
  1311 => (x"cd",x"c4",x"58",x"cc"),
  1312 => (x"78",x"c0",x"48",x"d4"),
  1313 => (x"de",x"dc",x"49",x"c1"),
  1314 => (x"1e",x"4f",x"26",x"87"),
  1315 => (x"d2",x"02",x"99",x"71"),
  1316 => (x"d8",x"f5",x"c1",x"87"),
  1317 => (x"f7",x"50",x"c0",x"48"),
  1318 => (x"ec",x"d1",x"c1",x"80"),
  1319 => (x"f4",x"f3",x"c1",x"40"),
  1320 => (x"c1",x"87",x"ce",x"78"),
  1321 => (x"c1",x"48",x"d4",x"f5"),
  1322 => (x"fc",x"78",x"ec",x"f3"),
  1323 => (x"e3",x"d1",x"c1",x"80"),
  1324 => (x"0e",x"4f",x"26",x"78"),
  1325 => (x"5d",x"5c",x"5b",x"5e"),
  1326 => (x"c3",x"86",x"f4",x"0e"),
  1327 => (x"c0",x"4d",x"d0",x"ff"),
  1328 => (x"48",x"a6",x"c8",x"4c"),
  1329 => (x"7e",x"75",x"78",x"c0"),
  1330 => (x"bf",x"d4",x"cd",x"c4"),
  1331 => (x"06",x"a8",x"c0",x"48"),
  1332 => (x"c8",x"87",x"c0",x"c1"),
  1333 => (x"7e",x"75",x"5c",x"a6"),
  1334 => (x"48",x"d0",x"ff",x"c3"),
  1335 => (x"f2",x"c0",x"02",x"98"),
  1336 => (x"4d",x"66",x"c4",x"87"),
  1337 => (x"1e",x"de",x"c5",x"c1"),
  1338 => (x"c4",x"02",x"66",x"cc"),
  1339 => (x"c2",x"4c",x"c0",x"87"),
  1340 => (x"74",x"4c",x"c1",x"87"),
  1341 => (x"87",x"f7",x"e0",x"49"),
  1342 => (x"7e",x"70",x"86",x"c4"),
  1343 => (x"66",x"c8",x"85",x"c1"),
  1344 => (x"cc",x"80",x"c1",x"48"),
  1345 => (x"cd",x"c4",x"58",x"a6"),
  1346 => (x"03",x"ad",x"bf",x"d4"),
  1347 => (x"05",x"6e",x"87",x"c5"),
  1348 => (x"6e",x"87",x"d1",x"ff"),
  1349 => (x"75",x"4c",x"c0",x"4d"),
  1350 => (x"dd",x"c3",x"02",x"9d"),
  1351 => (x"de",x"c5",x"c1",x"87"),
  1352 => (x"02",x"66",x"cc",x"1e"),
  1353 => (x"a6",x"c8",x"87",x"c7"),
  1354 => (x"c5",x"78",x"c0",x"48"),
  1355 => (x"48",x"a6",x"c8",x"87"),
  1356 => (x"66",x"c8",x"78",x"c1"),
  1357 => (x"f6",x"df",x"ff",x"49"),
  1358 => (x"70",x"86",x"c4",x"87"),
  1359 => (x"02",x"98",x"48",x"7e"),
  1360 => (x"49",x"87",x"e4",x"c2"),
  1361 => (x"69",x"97",x"81",x"cb"),
  1362 => (x"02",x"99",x"d0",x"49"),
  1363 => (x"74",x"87",x"d4",x"c1"),
  1364 => (x"c1",x"91",x"cc",x"49"),
  1365 => (x"c1",x"81",x"fc",x"f3"),
  1366 => (x"c8",x"79",x"fb",x"d0"),
  1367 => (x"51",x"ff",x"c3",x"81"),
  1368 => (x"91",x"de",x"49",x"74"),
  1369 => (x"4d",x"e8",x"cd",x"c4"),
  1370 => (x"c1",x"c2",x"85",x"71"),
  1371 => (x"a5",x"c1",x"7d",x"97"),
  1372 => (x"51",x"e0",x"c0",x"49"),
  1373 => (x"97",x"e0",x"c7",x"c4"),
  1374 => (x"87",x"d2",x"02",x"bf"),
  1375 => (x"a5",x"c2",x"84",x"c1"),
  1376 => (x"e0",x"c7",x"c4",x"4b"),
  1377 => (x"fe",x"49",x"db",x"4a"),
  1378 => (x"c1",x"87",x"f7",x"ec"),
  1379 => (x"a5",x"cd",x"87",x"d9"),
  1380 => (x"c1",x"51",x"c0",x"49"),
  1381 => (x"4b",x"a5",x"c2",x"84"),
  1382 => (x"49",x"cb",x"4a",x"6e"),
  1383 => (x"87",x"e2",x"ec",x"fe"),
  1384 => (x"74",x"87",x"c4",x"c1"),
  1385 => (x"c1",x"91",x"cc",x"49"),
  1386 => (x"c1",x"81",x"fc",x"f3"),
  1387 => (x"c4",x"79",x"ed",x"ce"),
  1388 => (x"bf",x"97",x"e0",x"c7"),
  1389 => (x"74",x"87",x"d8",x"02"),
  1390 => (x"c1",x"91",x"de",x"49"),
  1391 => (x"e8",x"cd",x"c4",x"84"),
  1392 => (x"c4",x"83",x"71",x"4b"),
  1393 => (x"dd",x"4a",x"e0",x"c7"),
  1394 => (x"f5",x"eb",x"fe",x"49"),
  1395 => (x"74",x"87",x"d8",x"87"),
  1396 => (x"c4",x"93",x"de",x"4b"),
  1397 => (x"cb",x"83",x"e8",x"cd"),
  1398 => (x"51",x"c0",x"49",x"a3"),
  1399 => (x"6e",x"73",x"84",x"c1"),
  1400 => (x"fe",x"49",x"cb",x"4a"),
  1401 => (x"c8",x"87",x"db",x"eb"),
  1402 => (x"80",x"c1",x"48",x"66"),
  1403 => (x"c7",x"58",x"a6",x"cc"),
  1404 => (x"c5",x"c0",x"03",x"ac"),
  1405 => (x"fc",x"05",x"6e",x"87"),
  1406 => (x"48",x"74",x"87",x"e3"),
  1407 => (x"4d",x"26",x"8e",x"f4"),
  1408 => (x"4b",x"26",x"4c",x"26"),
  1409 => (x"73",x"1e",x"4f",x"26"),
  1410 => (x"49",x"4b",x"71",x"1e"),
  1411 => (x"f3",x"c1",x"91",x"cc"),
  1412 => (x"a1",x"c8",x"81",x"fc"),
  1413 => (x"e0",x"f3",x"c1",x"4a"),
  1414 => (x"c9",x"50",x"12",x"48"),
  1415 => (x"c8",x"c1",x"4a",x"a1"),
  1416 => (x"50",x"12",x"48",x"c4"),
  1417 => (x"f3",x"c1",x"81",x"ca"),
  1418 => (x"50",x"11",x"48",x"e4"),
  1419 => (x"97",x"e4",x"f3",x"c1"),
  1420 => (x"c0",x"1e",x"49",x"bf"),
  1421 => (x"df",x"cc",x"c2",x"49"),
  1422 => (x"c8",x"cc",x"c4",x"87"),
  1423 => (x"c1",x"78",x"de",x"48"),
  1424 => (x"87",x"e3",x"d5",x"49"),
  1425 => (x"4b",x"26",x"8e",x"fc"),
  1426 => (x"5e",x"0e",x"4f",x"26"),
  1427 => (x"0e",x"5d",x"5c",x"5b"),
  1428 => (x"4d",x"71",x"86",x"f4"),
  1429 => (x"c1",x"91",x"cc",x"49"),
  1430 => (x"c8",x"81",x"fc",x"f3"),
  1431 => (x"a1",x"ca",x"4a",x"a1"),
  1432 => (x"48",x"a6",x"c4",x"7e"),
  1433 => (x"bf",x"e4",x"d1",x"c4"),
  1434 => (x"bf",x"97",x"6e",x"78"),
  1435 => (x"4c",x"66",x"c4",x"4b"),
  1436 => (x"48",x"12",x"2c",x"73"),
  1437 => (x"70",x"58",x"a6",x"cc"),
  1438 => (x"c9",x"84",x"c1",x"9c"),
  1439 => (x"49",x"69",x"97",x"81"),
  1440 => (x"c2",x"04",x"ac",x"b7"),
  1441 => (x"6e",x"4c",x"c0",x"87"),
  1442 => (x"c8",x"4a",x"bf",x"97"),
  1443 => (x"31",x"72",x"49",x"66"),
  1444 => (x"66",x"c4",x"b9",x"ff"),
  1445 => (x"72",x"48",x"74",x"99"),
  1446 => (x"48",x"4a",x"70",x"30"),
  1447 => (x"d1",x"c4",x"b0",x"71"),
  1448 => (x"f9",x"c1",x"58",x"e8"),
  1449 => (x"49",x"c0",x"87",x"f1"),
  1450 => (x"75",x"87",x"fc",x"d3"),
  1451 => (x"e7",x"fb",x"c0",x"49"),
  1452 => (x"26",x"8e",x"f4",x"87"),
  1453 => (x"26",x"4c",x"26",x"4d"),
  1454 => (x"1e",x"4f",x"26",x"4b"),
  1455 => (x"4b",x"71",x"1e",x"73"),
  1456 => (x"02",x"4a",x"a3",x"c6"),
  1457 => (x"8a",x"c1",x"87",x"db"),
  1458 => (x"8a",x"87",x"d6",x"02"),
  1459 => (x"87",x"da",x"c1",x"02"),
  1460 => (x"fc",x"c0",x"02",x"8a"),
  1461 => (x"c0",x"02",x"8a",x"87"),
  1462 => (x"02",x"8a",x"87",x"e1"),
  1463 => (x"db",x"c1",x"87",x"cb"),
  1464 => (x"f6",x"49",x"c7",x"87"),
  1465 => (x"de",x"c1",x"87",x"c6"),
  1466 => (x"d4",x"cd",x"c4",x"87"),
  1467 => (x"cb",x"c1",x"02",x"bf"),
  1468 => (x"88",x"c1",x"48",x"87"),
  1469 => (x"58",x"d8",x"cd",x"c4"),
  1470 => (x"c4",x"87",x"c1",x"c1"),
  1471 => (x"02",x"bf",x"d8",x"cd"),
  1472 => (x"c4",x"87",x"f9",x"c0"),
  1473 => (x"48",x"bf",x"d4",x"cd"),
  1474 => (x"cd",x"c4",x"80",x"c1"),
  1475 => (x"eb",x"c0",x"58",x"d8"),
  1476 => (x"d4",x"cd",x"c4",x"87"),
  1477 => (x"89",x"c6",x"49",x"bf"),
  1478 => (x"59",x"d8",x"cd",x"c4"),
  1479 => (x"03",x"a9",x"b7",x"c0"),
  1480 => (x"cd",x"c4",x"87",x"da"),
  1481 => (x"78",x"c0",x"48",x"d4"),
  1482 => (x"cd",x"c4",x"87",x"d2"),
  1483 => (x"cb",x"02",x"bf",x"d8"),
  1484 => (x"d4",x"cd",x"c4",x"87"),
  1485 => (x"80",x"c6",x"48",x"bf"),
  1486 => (x"58",x"d8",x"cd",x"c4"),
  1487 => (x"e6",x"d1",x"49",x"c0"),
  1488 => (x"c0",x"49",x"73",x"87"),
  1489 => (x"26",x"87",x"d1",x"f9"),
  1490 => (x"0e",x"4f",x"26",x"4b"),
  1491 => (x"5d",x"5c",x"5b",x"5e"),
  1492 => (x"86",x"d4",x"ff",x"0e"),
  1493 => (x"c8",x"59",x"a6",x"dc"),
  1494 => (x"78",x"c0",x"48",x"a6"),
  1495 => (x"c0",x"c1",x"80",x"c4"),
  1496 => (x"80",x"c4",x"78",x"66"),
  1497 => (x"80",x"c4",x"78",x"c1"),
  1498 => (x"cd",x"c4",x"78",x"c1"),
  1499 => (x"78",x"c1",x"48",x"d8"),
  1500 => (x"bf",x"c8",x"cc",x"c4"),
  1501 => (x"05",x"a8",x"de",x"48"),
  1502 => (x"f6",x"f4",x"87",x"c9"),
  1503 => (x"58",x"a6",x"cc",x"87"),
  1504 => (x"c1",x"87",x"df",x"cf"),
  1505 => (x"e4",x"87",x"ec",x"f7"),
  1506 => (x"f7",x"c1",x"87",x"e8"),
  1507 => (x"4c",x"70",x"87",x"c2"),
  1508 => (x"02",x"ac",x"fb",x"c0"),
  1509 => (x"d8",x"87",x"f0",x"c1"),
  1510 => (x"e2",x"c1",x"05",x"66"),
  1511 => (x"66",x"fc",x"c0",x"87"),
  1512 => (x"6a",x"82",x"c4",x"4a"),
  1513 => (x"d8",x"ee",x"c1",x"7e"),
  1514 => (x"20",x"49",x"6e",x"48"),
  1515 => (x"10",x"41",x"20",x"41"),
  1516 => (x"66",x"fc",x"c0",x"51"),
  1517 => (x"c6",x"d8",x"c1",x"48"),
  1518 => (x"c7",x"49",x"6a",x"78"),
  1519 => (x"c0",x"51",x"74",x"81"),
  1520 => (x"c8",x"49",x"66",x"fc"),
  1521 => (x"c0",x"51",x"c1",x"81"),
  1522 => (x"c9",x"49",x"66",x"fc"),
  1523 => (x"c0",x"51",x"c0",x"81"),
  1524 => (x"ca",x"49",x"66",x"fc"),
  1525 => (x"c1",x"51",x"c0",x"81"),
  1526 => (x"6a",x"1e",x"d8",x"1e"),
  1527 => (x"e3",x"81",x"c8",x"49"),
  1528 => (x"86",x"c8",x"87",x"e5"),
  1529 => (x"48",x"66",x"c0",x"c1"),
  1530 => (x"c7",x"01",x"a8",x"c0"),
  1531 => (x"48",x"a6",x"c8",x"87"),
  1532 => (x"87",x"ce",x"78",x"c1"),
  1533 => (x"48",x"66",x"c0",x"c1"),
  1534 => (x"a6",x"d0",x"88",x"c1"),
  1535 => (x"e2",x"87",x"c3",x"58"),
  1536 => (x"a6",x"d0",x"87",x"f0"),
  1537 => (x"74",x"78",x"c2",x"48"),
  1538 => (x"d1",x"cd",x"02",x"9c"),
  1539 => (x"48",x"66",x"c8",x"87"),
  1540 => (x"a8",x"66",x"c4",x"c1"),
  1541 => (x"87",x"c6",x"cd",x"03"),
  1542 => (x"c0",x"48",x"a6",x"dc"),
  1543 => (x"f4",x"c1",x"7e",x"78"),
  1544 => (x"4c",x"70",x"87",x"ee"),
  1545 => (x"05",x"ac",x"d0",x"c1"),
  1546 => (x"c4",x"87",x"d9",x"c2"),
  1547 => (x"78",x"6e",x"48",x"a6"),
  1548 => (x"70",x"87",x"c1",x"e4"),
  1549 => (x"d7",x"f4",x"c1",x"7e"),
  1550 => (x"c0",x"4c",x"70",x"87"),
  1551 => (x"c1",x"05",x"ac",x"ec"),
  1552 => (x"66",x"c8",x"87",x"ed"),
  1553 => (x"c0",x"91",x"cc",x"49"),
  1554 => (x"c4",x"81",x"66",x"fc"),
  1555 => (x"4d",x"6a",x"4a",x"a1"),
  1556 => (x"6e",x"4a",x"a1",x"c8"),
  1557 => (x"ec",x"d1",x"c1",x"52"),
  1558 => (x"f3",x"f3",x"c1",x"79"),
  1559 => (x"9c",x"4c",x"70",x"87"),
  1560 => (x"c0",x"87",x"d9",x"02"),
  1561 => (x"d3",x"02",x"ac",x"fb"),
  1562 => (x"c1",x"55",x"74",x"87"),
  1563 => (x"70",x"87",x"e1",x"f3"),
  1564 => (x"c7",x"02",x"9c",x"4c"),
  1565 => (x"ac",x"fb",x"c0",x"87"),
  1566 => (x"87",x"ed",x"ff",x"05"),
  1567 => (x"c2",x"55",x"e0",x"c0"),
  1568 => (x"97",x"c0",x"55",x"c1"),
  1569 => (x"48",x"66",x"d8",x"7d"),
  1570 => (x"05",x"a8",x"66",x"c4"),
  1571 => (x"66",x"c8",x"87",x"db"),
  1572 => (x"a8",x"66",x"cc",x"48"),
  1573 => (x"c8",x"87",x"ca",x"04"),
  1574 => (x"80",x"c1",x"48",x"66"),
  1575 => (x"c8",x"58",x"a6",x"cc"),
  1576 => (x"48",x"66",x"cc",x"87"),
  1577 => (x"a6",x"d0",x"88",x"c1"),
  1578 => (x"e3",x"f2",x"c1",x"58"),
  1579 => (x"c1",x"4c",x"70",x"87"),
  1580 => (x"c8",x"05",x"ac",x"d0"),
  1581 => (x"48",x"66",x"d4",x"87"),
  1582 => (x"a6",x"d8",x"80",x"c1"),
  1583 => (x"ac",x"d0",x"c1",x"58"),
  1584 => (x"87",x"e7",x"fd",x"02"),
  1585 => (x"66",x"d8",x"48",x"6e"),
  1586 => (x"e3",x"c9",x"05",x"a8"),
  1587 => (x"a6",x"e0",x"c0",x"87"),
  1588 => (x"74",x"78",x"c0",x"48"),
  1589 => (x"88",x"fb",x"c0",x"48"),
  1590 => (x"70",x"58",x"a6",x"c8"),
  1591 => (x"e4",x"c9",x"02",x"98"),
  1592 => (x"88",x"cb",x"48",x"87"),
  1593 => (x"70",x"58",x"a6",x"c8"),
  1594 => (x"d1",x"c1",x"02",x"98"),
  1595 => (x"88",x"c9",x"48",x"87"),
  1596 => (x"70",x"58",x"a6",x"c8"),
  1597 => (x"c1",x"c4",x"02",x"98"),
  1598 => (x"88",x"c4",x"48",x"87"),
  1599 => (x"70",x"58",x"a6",x"c8"),
  1600 => (x"87",x"cf",x"02",x"98"),
  1601 => (x"c8",x"88",x"c1",x"48"),
  1602 => (x"98",x"70",x"58",x"a6"),
  1603 => (x"87",x"ea",x"c3",x"02"),
  1604 => (x"dc",x"87",x"d4",x"c8"),
  1605 => (x"f0",x"c0",x"48",x"a6"),
  1606 => (x"f3",x"f0",x"c1",x"78"),
  1607 => (x"c0",x"4c",x"70",x"87"),
  1608 => (x"c0",x"02",x"ac",x"ec"),
  1609 => (x"e0",x"c0",x"87",x"c4"),
  1610 => (x"ec",x"c0",x"5c",x"a6"),
  1611 => (x"cd",x"c0",x"02",x"ac"),
  1612 => (x"db",x"f0",x"c1",x"87"),
  1613 => (x"c0",x"4c",x"70",x"87"),
  1614 => (x"ff",x"05",x"ac",x"ec"),
  1615 => (x"ec",x"c0",x"87",x"f3"),
  1616 => (x"c4",x"c0",x"02",x"ac"),
  1617 => (x"c7",x"f0",x"c1",x"87"),
  1618 => (x"ca",x"1e",x"c0",x"87"),
  1619 => (x"49",x"66",x"d0",x"1e"),
  1620 => (x"c4",x"c1",x"91",x"cc"),
  1621 => (x"80",x"71",x"48",x"66"),
  1622 => (x"c8",x"58",x"a6",x"cc"),
  1623 => (x"80",x"c4",x"48",x"66"),
  1624 => (x"cc",x"58",x"a6",x"d0"),
  1625 => (x"ff",x"49",x"bf",x"66"),
  1626 => (x"c1",x"87",x"dc",x"dd"),
  1627 => (x"d4",x"1e",x"de",x"1e"),
  1628 => (x"ff",x"49",x"bf",x"66"),
  1629 => (x"d0",x"87",x"d0",x"dd"),
  1630 => (x"48",x"49",x"70",x"86"),
  1631 => (x"c0",x"88",x"08",x"c0"),
  1632 => (x"c0",x"58",x"a6",x"e8"),
  1633 => (x"ee",x"c0",x"06",x"a8"),
  1634 => (x"66",x"e4",x"c0",x"87"),
  1635 => (x"03",x"a8",x"dd",x"48"),
  1636 => (x"c4",x"87",x"e4",x"c0"),
  1637 => (x"c0",x"49",x"bf",x"66"),
  1638 => (x"c0",x"81",x"66",x"e4"),
  1639 => (x"e4",x"c0",x"51",x"e0"),
  1640 => (x"81",x"c1",x"49",x"66"),
  1641 => (x"81",x"bf",x"66",x"c4"),
  1642 => (x"c0",x"51",x"c1",x"c2"),
  1643 => (x"c2",x"49",x"66",x"e4"),
  1644 => (x"bf",x"66",x"c4",x"81"),
  1645 => (x"6e",x"51",x"c0",x"81"),
  1646 => (x"c6",x"d8",x"c1",x"48"),
  1647 => (x"c8",x"49",x"6e",x"78"),
  1648 => (x"51",x"66",x"d0",x"81"),
  1649 => (x"81",x"c9",x"49",x"6e"),
  1650 => (x"6e",x"51",x"66",x"d4"),
  1651 => (x"dc",x"81",x"ca",x"49"),
  1652 => (x"66",x"d0",x"51",x"66"),
  1653 => (x"d4",x"80",x"c1",x"48"),
  1654 => (x"66",x"c8",x"58",x"a6"),
  1655 => (x"a8",x"66",x"cc",x"48"),
  1656 => (x"87",x"cb",x"c0",x"04"),
  1657 => (x"c1",x"48",x"66",x"c8"),
  1658 => (x"58",x"a6",x"cc",x"80"),
  1659 => (x"cc",x"87",x"d6",x"c5"),
  1660 => (x"88",x"c1",x"48",x"66"),
  1661 => (x"c5",x"58",x"a6",x"d0"),
  1662 => (x"dc",x"ff",x"87",x"cb"),
  1663 => (x"e8",x"c0",x"87",x"f6"),
  1664 => (x"dc",x"ff",x"58",x"a6"),
  1665 => (x"e0",x"c0",x"87",x"ee"),
  1666 => (x"ec",x"c0",x"58",x"a6"),
  1667 => (x"ca",x"c0",x"05",x"a8"),
  1668 => (x"48",x"a6",x"dc",x"87"),
  1669 => (x"78",x"66",x"e4",x"c0"),
  1670 => (x"c1",x"87",x"c4",x"c0"),
  1671 => (x"c8",x"87",x"f1",x"ec"),
  1672 => (x"91",x"cc",x"49",x"66"),
  1673 => (x"48",x"66",x"fc",x"c0"),
  1674 => (x"a6",x"c8",x"80",x"71"),
  1675 => (x"4a",x"66",x"c4",x"58"),
  1676 => (x"66",x"c4",x"82",x"c8"),
  1677 => (x"c0",x"81",x"ca",x"49"),
  1678 => (x"dc",x"51",x"66",x"e4"),
  1679 => (x"81",x"c1",x"49",x"66"),
  1680 => (x"89",x"66",x"e4",x"c0"),
  1681 => (x"30",x"71",x"48",x"c1"),
  1682 => (x"89",x"c1",x"49",x"70"),
  1683 => (x"c4",x"7a",x"97",x"71"),
  1684 => (x"49",x"bf",x"e4",x"d1"),
  1685 => (x"29",x"66",x"e4",x"c0"),
  1686 => (x"48",x"4a",x"6a",x"97"),
  1687 => (x"ec",x"c0",x"98",x"71"),
  1688 => (x"66",x"c4",x"58",x"a6"),
  1689 => (x"69",x"81",x"c4",x"49"),
  1690 => (x"48",x"66",x"d8",x"4d"),
  1691 => (x"c0",x"02",x"a8",x"6e"),
  1692 => (x"7e",x"c0",x"87",x"c5"),
  1693 => (x"c1",x"87",x"c2",x"c0"),
  1694 => (x"c0",x"1e",x"6e",x"7e"),
  1695 => (x"49",x"75",x"1e",x"e0"),
  1696 => (x"87",x"c3",x"d9",x"ff"),
  1697 => (x"4c",x"70",x"86",x"c8"),
  1698 => (x"06",x"ac",x"b7",x"c0"),
  1699 => (x"74",x"87",x"d0",x"c1"),
  1700 => (x"49",x"e0",x"c0",x"85"),
  1701 => (x"4b",x"75",x"89",x"74"),
  1702 => (x"4a",x"e4",x"ee",x"c1"),
  1703 => (x"e1",x"d8",x"fe",x"71"),
  1704 => (x"75",x"85",x"c2",x"87"),
  1705 => (x"66",x"e0",x"c0",x"7e"),
  1706 => (x"c0",x"80",x"c1",x"48"),
  1707 => (x"c0",x"58",x"a6",x"e4"),
  1708 => (x"c1",x"49",x"66",x"e8"),
  1709 => (x"02",x"a9",x"70",x"81"),
  1710 => (x"c0",x"87",x"c5",x"c0"),
  1711 => (x"87",x"c2",x"c0",x"4d"),
  1712 => (x"1e",x"75",x"4d",x"c1"),
  1713 => (x"c0",x"49",x"a4",x"c2"),
  1714 => (x"88",x"71",x"48",x"e0"),
  1715 => (x"c8",x"1e",x"49",x"70"),
  1716 => (x"d7",x"ff",x"49",x"66"),
  1717 => (x"86",x"c8",x"87",x"f1"),
  1718 => (x"01",x"a8",x"b7",x"c0"),
  1719 => (x"c0",x"87",x"c6",x"ff"),
  1720 => (x"c0",x"02",x"66",x"e0"),
  1721 => (x"66",x"c4",x"87",x"d3"),
  1722 => (x"c0",x"81",x"c9",x"49"),
  1723 => (x"c4",x"51",x"66",x"e0"),
  1724 => (x"d9",x"c1",x"48",x"66"),
  1725 => (x"ce",x"c0",x"78",x"ca"),
  1726 => (x"49",x"66",x"c4",x"87"),
  1727 => (x"51",x"c2",x"81",x"c9"),
  1728 => (x"c3",x"48",x"66",x"c4"),
  1729 => (x"c8",x"78",x"d0",x"dd"),
  1730 => (x"66",x"cc",x"48",x"66"),
  1731 => (x"cb",x"c0",x"04",x"a8"),
  1732 => (x"48",x"66",x"c8",x"87"),
  1733 => (x"a6",x"cc",x"80",x"c1"),
  1734 => (x"87",x"e9",x"c0",x"58"),
  1735 => (x"c1",x"48",x"66",x"cc"),
  1736 => (x"58",x"a6",x"d0",x"88"),
  1737 => (x"ff",x"87",x"de",x"c0"),
  1738 => (x"70",x"87",x"c7",x"d6"),
  1739 => (x"87",x"d5",x"c0",x"4c"),
  1740 => (x"05",x"ac",x"c6",x"c1"),
  1741 => (x"d0",x"87",x"c8",x"c0"),
  1742 => (x"80",x"c1",x"48",x"66"),
  1743 => (x"ff",x"58",x"a6",x"d4"),
  1744 => (x"70",x"87",x"ef",x"d5"),
  1745 => (x"48",x"66",x"d4",x"4c"),
  1746 => (x"a6",x"d8",x"80",x"c1"),
  1747 => (x"02",x"9c",x"74",x"58"),
  1748 => (x"c8",x"87",x"cb",x"c0"),
  1749 => (x"c4",x"c1",x"48",x"66"),
  1750 => (x"f2",x"04",x"a8",x"66"),
  1751 => (x"d5",x"ff",x"87",x"fa"),
  1752 => (x"66",x"c8",x"87",x"c7"),
  1753 => (x"03",x"a8",x"c7",x"48"),
  1754 => (x"c8",x"87",x"e1",x"c0"),
  1755 => (x"cd",x"c4",x"4c",x"66"),
  1756 => (x"78",x"c0",x"48",x"d8"),
  1757 => (x"91",x"cc",x"49",x"74"),
  1758 => (x"81",x"66",x"fc",x"c0"),
  1759 => (x"6a",x"4a",x"a1",x"c4"),
  1760 => (x"79",x"52",x"c0",x"4a"),
  1761 => (x"ac",x"c7",x"84",x"c1"),
  1762 => (x"87",x"e2",x"ff",x"04"),
  1763 => (x"26",x"8e",x"d4",x"ff"),
  1764 => (x"26",x"4c",x"26",x"4d"),
  1765 => (x"00",x"4f",x"26",x"4b"),
  1766 => (x"64",x"61",x"6f",x"4c"),
  1767 => (x"20",x"2e",x"2a",x"20"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"1e",x"00",x"20",x"3a"),
  1770 => (x"4b",x"71",x"1e",x"73"),
  1771 => (x"87",x"c6",x"02",x"9b"),
  1772 => (x"48",x"d4",x"cd",x"c4"),
  1773 => (x"1e",x"c7",x"78",x"c0"),
  1774 => (x"bf",x"d4",x"cd",x"c4"),
  1775 => (x"fc",x"f3",x"c1",x"1e"),
  1776 => (x"c8",x"cc",x"c4",x"1e"),
  1777 => (x"c2",x"ee",x"49",x"bf"),
  1778 => (x"c4",x"86",x"cc",x"87"),
  1779 => (x"49",x"bf",x"c8",x"cc"),
  1780 => (x"73",x"87",x"f8",x"e2"),
  1781 => (x"87",x"c8",x"02",x"9b"),
  1782 => (x"49",x"fc",x"f3",x"c1"),
  1783 => (x"87",x"c6",x"e8",x"c0"),
  1784 => (x"4f",x"26",x"4b",x"26"),
  1785 => (x"fc",x"1e",x"73",x"1e"),
  1786 => (x"4b",x"ff",x"c3",x"86"),
  1787 => (x"fc",x"4a",x"d4",x"ff"),
  1788 => (x"98",x"c1",x"48",x"bf"),
  1789 => (x"98",x"48",x"7e",x"70"),
  1790 => (x"87",x"fb",x"c0",x"02"),
  1791 => (x"c1",x"48",x"d0",x"ff"),
  1792 => (x"d2",x"c2",x"78",x"c1"),
  1793 => (x"c3",x"7a",x"73",x"7a"),
  1794 => (x"48",x"49",x"d1",x"ff"),
  1795 => (x"50",x"6a",x"80",x"ff"),
  1796 => (x"51",x"6a",x"7a",x"73"),
  1797 => (x"80",x"c1",x"7a",x"73"),
  1798 => (x"7a",x"73",x"50",x"6a"),
  1799 => (x"7a",x"73",x"50",x"6a"),
  1800 => (x"7a",x"73",x"49",x"6a"),
  1801 => (x"7a",x"73",x"50",x"6a"),
  1802 => (x"ff",x"c3",x"50",x"6a"),
  1803 => (x"ff",x"59",x"97",x"da"),
  1804 => (x"c0",x"c1",x"48",x"d0"),
  1805 => (x"c3",x"87",x"d7",x"78"),
  1806 => (x"48",x"49",x"d1",x"ff"),
  1807 => (x"50",x"c0",x"80",x"ff"),
  1808 => (x"c0",x"80",x"c1",x"51"),
  1809 => (x"c1",x"50",x"d9",x"50"),
  1810 => (x"50",x"e2",x"c0",x"50"),
  1811 => (x"ff",x"c3",x"50",x"c3"),
  1812 => (x"50",x"c0",x"48",x"d7"),
  1813 => (x"8e",x"fc",x"80",x"f8"),
  1814 => (x"4f",x"26",x"4b",x"26"),
  1815 => (x"87",x"d0",x"cc",x"1e"),
  1816 => (x"c2",x"fd",x"49",x"c1"),
  1817 => (x"d1",x"dc",x"fe",x"87"),
  1818 => (x"02",x"98",x"70",x"87"),
  1819 => (x"e5",x"fe",x"87",x"cd"),
  1820 => (x"98",x"70",x"87",x"dd"),
  1821 => (x"c1",x"87",x"c4",x"02"),
  1822 => (x"c0",x"87",x"c2",x"4a"),
  1823 => (x"05",x"9a",x"72",x"4a"),
  1824 => (x"1e",x"c0",x"87",x"ce"),
  1825 => (x"49",x"f0",x"f2",x"c1"),
  1826 => (x"87",x"e5",x"f2",x"c0"),
  1827 => (x"87",x"fe",x"86",x"c4"),
  1828 => (x"f2",x"c1",x"1e",x"c0"),
  1829 => (x"f2",x"c0",x"49",x"fc"),
  1830 => (x"1e",x"c0",x"87",x"d7"),
  1831 => (x"87",x"c2",x"f9",x"c1"),
  1832 => (x"f2",x"c0",x"49",x"70"),
  1833 => (x"d2",x"c3",x"87",x"cb"),
  1834 => (x"26",x"8e",x"f8",x"87"),
  1835 => (x"00",x"00",x"00",x"4f"),
  1836 => (x"66",x"20",x"44",x"53"),
  1837 => (x"65",x"6c",x"69",x"61"),
  1838 => (x"00",x"00",x"2e",x"64"),
  1839 => (x"74",x"6f",x"6f",x"42"),
  1840 => (x"2e",x"67",x"6e",x"69"),
  1841 => (x"1e",x"00",x"2e",x"2e"),
  1842 => (x"48",x"d4",x"cd",x"c4"),
  1843 => (x"cc",x"c4",x"78",x"c0"),
  1844 => (x"78",x"c0",x"48",x"c8"),
  1845 => (x"c1",x"87",x"c5",x"fe"),
  1846 => (x"c0",x"87",x"e4",x"fb"),
  1847 => (x"00",x"4f",x"26",x"48"),
  1848 => (x"00",x"00",x"00",x"00"),
  1849 => (x"00",x"00",x"00",x"00"),
  1850 => (x"00",x"00",x"00",x"01"),
  1851 => (x"78",x"45",x"20",x"80"),
  1852 => (x"00",x"00",x"74",x"69"),
  1853 => (x"61",x"42",x"20",x"80"),
  1854 => (x"00",x"00",x"6b",x"63"),
  1855 => (x"00",x"00",x"13",x"ad"),
  1856 => (x"00",x"00",x"43",x"68"),
  1857 => (x"00",x"00",x"00",x"00"),
  1858 => (x"00",x"00",x"13",x"ad"),
  1859 => (x"00",x"00",x"43",x"86"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"13",x"ad"),
  1862 => (x"00",x"00",x"43",x"a4"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"13",x"ad"),
  1865 => (x"00",x"00",x"43",x"c2"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"13",x"ad"),
  1868 => (x"00",x"00",x"43",x"e0"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"13",x"ad"),
  1871 => (x"00",x"00",x"43",x"fe"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"13",x"ad"),
  1874 => (x"00",x"00",x"44",x"1c"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"14",x"6c"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"16",x"bb"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"48",x"f0",x"fe",x"1e"),
  1883 => (x"09",x"cd",x"78",x"c0"),
  1884 => (x"4f",x"26",x"09",x"79"),
  1885 => (x"bf",x"f0",x"fe",x"1e"),
  1886 => (x"1e",x"4f",x"26",x"48"),
  1887 => (x"c1",x"48",x"f0",x"fe"),
  1888 => (x"1e",x"4f",x"26",x"78"),
  1889 => (x"c0",x"48",x"f0",x"fe"),
  1890 => (x"1e",x"4f",x"26",x"78"),
  1891 => (x"97",x"c0",x"4a",x"71"),
  1892 => (x"49",x"a2",x"c1",x"7a"),
  1893 => (x"a2",x"ca",x"51",x"c0"),
  1894 => (x"cb",x"51",x"c0",x"49"),
  1895 => (x"51",x"c0",x"49",x"a2"),
  1896 => (x"5e",x"0e",x"4f",x"26"),
  1897 => (x"f0",x"0e",x"5c",x"5b"),
  1898 => (x"ca",x"4c",x"71",x"86"),
  1899 => (x"69",x"97",x"49",x"a4"),
  1900 => (x"4b",x"a4",x"cb",x"7e"),
  1901 => (x"c8",x"48",x"6b",x"97"),
  1902 => (x"80",x"c1",x"58",x"a6"),
  1903 => (x"c7",x"58",x"a6",x"cc"),
  1904 => (x"58",x"a6",x"d0",x"98"),
  1905 => (x"66",x"cc",x"48",x"6e"),
  1906 => (x"87",x"db",x"05",x"a8"),
  1907 => (x"97",x"7e",x"69",x"97"),
  1908 => (x"a6",x"c8",x"48",x"6b"),
  1909 => (x"cc",x"80",x"c1",x"58"),
  1910 => (x"98",x"c7",x"58",x"a6"),
  1911 => (x"6e",x"58",x"a6",x"d0"),
  1912 => (x"a8",x"66",x"cc",x"48"),
  1913 => (x"fe",x"87",x"e5",x"02"),
  1914 => (x"a4",x"cc",x"87",x"d9"),
  1915 => (x"49",x"6b",x"97",x"4a"),
  1916 => (x"dc",x"49",x"a1",x"72"),
  1917 => (x"6b",x"97",x"51",x"66"),
  1918 => (x"c1",x"48",x"6e",x"7e"),
  1919 => (x"58",x"a6",x"c8",x"80"),
  1920 => (x"a6",x"cc",x"98",x"c7"),
  1921 => (x"7b",x"97",x"70",x"58"),
  1922 => (x"fd",x"87",x"d1",x"c2"),
  1923 => (x"8e",x"f0",x"87",x"ed"),
  1924 => (x"4b",x"26",x"4c",x"26"),
  1925 => (x"5e",x"0e",x"4f",x"26"),
  1926 => (x"0e",x"5d",x"5c",x"5b"),
  1927 => (x"4d",x"71",x"86",x"f4"),
  1928 => (x"c1",x"7e",x"6d",x"97"),
  1929 => (x"6c",x"97",x"4c",x"a5"),
  1930 => (x"58",x"a6",x"c8",x"48"),
  1931 => (x"66",x"c4",x"48",x"6e"),
  1932 => (x"87",x"c5",x"05",x"a8"),
  1933 => (x"e6",x"c0",x"48",x"ff"),
  1934 => (x"87",x"c7",x"fd",x"87"),
  1935 => (x"97",x"49",x"a5",x"c2"),
  1936 => (x"a3",x"71",x"4b",x"6c"),
  1937 => (x"4b",x"6b",x"97",x"4b"),
  1938 => (x"6e",x"7e",x"6c",x"97"),
  1939 => (x"c8",x"80",x"c1",x"48"),
  1940 => (x"98",x"c7",x"58",x"a6"),
  1941 => (x"70",x"58",x"a6",x"cc"),
  1942 => (x"de",x"fc",x"7c",x"97"),
  1943 => (x"f4",x"48",x"73",x"87"),
  1944 => (x"26",x"4d",x"26",x"8e"),
  1945 => (x"26",x"4b",x"26",x"4c"),
  1946 => (x"5b",x"5e",x"0e",x"4f"),
  1947 => (x"86",x"f4",x"0e",x"5c"),
  1948 => (x"66",x"d8",x"4c",x"71"),
  1949 => (x"9a",x"ff",x"c3",x"4a"),
  1950 => (x"97",x"4b",x"a4",x"c2"),
  1951 => (x"a1",x"73",x"49",x"6c"),
  1952 => (x"97",x"51",x"72",x"49"),
  1953 => (x"48",x"6e",x"7e",x"6c"),
  1954 => (x"a6",x"c8",x"80",x"c1"),
  1955 => (x"cc",x"98",x"c7",x"58"),
  1956 => (x"54",x"70",x"58",x"a6"),
  1957 => (x"4c",x"26",x"8e",x"f4"),
  1958 => (x"4f",x"26",x"4b",x"26"),
  1959 => (x"f4",x"1e",x"73",x"1e"),
  1960 => (x"87",x"df",x"fb",x"86"),
  1961 => (x"49",x"4b",x"bf",x"e0"),
  1962 => (x"99",x"c0",x"e0",x"c0"),
  1963 => (x"73",x"87",x"cb",x"02"),
  1964 => (x"fc",x"d0",x"c4",x"1e"),
  1965 => (x"87",x"f1",x"fe",x"49"),
  1966 => (x"49",x"73",x"86",x"c4"),
  1967 => (x"02",x"99",x"c0",x"d0"),
  1968 => (x"c4",x"87",x"c0",x"c1"),
  1969 => (x"bf",x"97",x"c6",x"d1"),
  1970 => (x"c7",x"d1",x"c4",x"7e"),
  1971 => (x"c8",x"48",x"bf",x"97"),
  1972 => (x"48",x"6e",x"58",x"a6"),
  1973 => (x"02",x"a8",x"66",x"c4"),
  1974 => (x"c4",x"87",x"e8",x"c0"),
  1975 => (x"bf",x"97",x"c6",x"d1"),
  1976 => (x"c8",x"d1",x"c4",x"49"),
  1977 => (x"e0",x"48",x"11",x"81"),
  1978 => (x"d1",x"c4",x"78",x"08"),
  1979 => (x"7e",x"bf",x"97",x"c6"),
  1980 => (x"80",x"c1",x"48",x"6e"),
  1981 => (x"c7",x"58",x"a6",x"c8"),
  1982 => (x"58",x"a6",x"cc",x"98"),
  1983 => (x"48",x"c6",x"d1",x"c4"),
  1984 => (x"e4",x"50",x"66",x"c8"),
  1985 => (x"c0",x"49",x"4b",x"bf"),
  1986 => (x"02",x"99",x"c0",x"e0"),
  1987 => (x"1e",x"73",x"87",x"cb"),
  1988 => (x"49",x"d0",x"d1",x"c4"),
  1989 => (x"c4",x"87",x"d2",x"fd"),
  1990 => (x"d0",x"49",x"73",x"86"),
  1991 => (x"c1",x"02",x"99",x"c0"),
  1992 => (x"d1",x"c4",x"87",x"c0"),
  1993 => (x"7e",x"bf",x"97",x"da"),
  1994 => (x"97",x"db",x"d1",x"c4"),
  1995 => (x"a6",x"c8",x"48",x"bf"),
  1996 => (x"c4",x"48",x"6e",x"58"),
  1997 => (x"c0",x"02",x"a8",x"66"),
  1998 => (x"d1",x"c4",x"87",x"e8"),
  1999 => (x"49",x"bf",x"97",x"da"),
  2000 => (x"81",x"dc",x"d1",x"c4"),
  2001 => (x"08",x"e4",x"48",x"11"),
  2002 => (x"da",x"d1",x"c4",x"78"),
  2003 => (x"6e",x"7e",x"bf",x"97"),
  2004 => (x"c8",x"80",x"c1",x"48"),
  2005 => (x"98",x"c7",x"58",x"a6"),
  2006 => (x"c4",x"58",x"a6",x"cc"),
  2007 => (x"c8",x"48",x"da",x"d1"),
  2008 => (x"cf",x"f8",x"50",x"66"),
  2009 => (x"f8",x"7e",x"70",x"87"),
  2010 => (x"8e",x"f4",x"87",x"d1"),
  2011 => (x"4f",x"26",x"4b",x"26"),
  2012 => (x"fc",x"d0",x"c4",x"1e"),
  2013 => (x"87",x"d3",x"f8",x"49"),
  2014 => (x"49",x"d0",x"d1",x"c4"),
  2015 => (x"c1",x"87",x"cc",x"f8"),
  2016 => (x"f7",x"49",x"dc",x"fa"),
  2017 => (x"ef",x"c2",x"87",x"e2"),
  2018 => (x"1e",x"4f",x"26",x"87"),
  2019 => (x"d0",x"c4",x"1e",x"73"),
  2020 => (x"c1",x"fa",x"49",x"fc"),
  2021 => (x"c0",x"4a",x"70",x"87"),
  2022 => (x"c2",x"04",x"aa",x"b7"),
  2023 => (x"f0",x"c3",x"87",x"cc"),
  2024 => (x"87",x"c9",x"05",x"aa"),
  2025 => (x"48",x"f0",x"c0",x"c2"),
  2026 => (x"ed",x"c1",x"78",x"c1"),
  2027 => (x"aa",x"e0",x"c3",x"87"),
  2028 => (x"c2",x"87",x"c9",x"05"),
  2029 => (x"c1",x"48",x"f4",x"c0"),
  2030 => (x"87",x"de",x"c1",x"78"),
  2031 => (x"bf",x"f4",x"c0",x"c2"),
  2032 => (x"c2",x"87",x"c6",x"02"),
  2033 => (x"c2",x"4b",x"a2",x"c0"),
  2034 => (x"c2",x"4b",x"72",x"87"),
  2035 => (x"02",x"bf",x"f0",x"c0"),
  2036 => (x"73",x"87",x"e0",x"c0"),
  2037 => (x"29",x"b7",x"c4",x"49"),
  2038 => (x"cc",x"c2",x"c2",x"91"),
  2039 => (x"cf",x"4a",x"73",x"81"),
  2040 => (x"c1",x"92",x"c2",x"9a"),
  2041 => (x"70",x"30",x"72",x"48"),
  2042 => (x"72",x"ba",x"ff",x"4a"),
  2043 => (x"70",x"98",x"69",x"48"),
  2044 => (x"73",x"87",x"db",x"79"),
  2045 => (x"29",x"b7",x"c4",x"49"),
  2046 => (x"cc",x"c2",x"c2",x"91"),
  2047 => (x"cf",x"4a",x"73",x"81"),
  2048 => (x"c3",x"92",x"c2",x"9a"),
  2049 => (x"70",x"30",x"72",x"48"),
  2050 => (x"b0",x"69",x"48",x"4a"),
  2051 => (x"c0",x"c2",x"79",x"70"),
  2052 => (x"78",x"c0",x"48",x"f4"),
  2053 => (x"48",x"f0",x"c0",x"c2"),
  2054 => (x"d0",x"c4",x"78",x"c0"),
  2055 => (x"f5",x"f7",x"49",x"fc"),
  2056 => (x"c0",x"4a",x"70",x"87"),
  2057 => (x"fd",x"03",x"aa",x"b7"),
  2058 => (x"48",x"c0",x"87",x"f4"),
  2059 => (x"4f",x"26",x"4b",x"26"),
  2060 => (x"00",x"00",x"00",x"00"),
  2061 => (x"00",x"00",x"00",x"00"),
  2062 => (x"72",x"4a",x"c0",x"1e"),
  2063 => (x"c2",x"91",x"c4",x"49"),
  2064 => (x"c0",x"81",x"cc",x"c2"),
  2065 => (x"d0",x"82",x"c1",x"79"),
  2066 => (x"ee",x"04",x"aa",x"b7"),
  2067 => (x"0e",x"4f",x"26",x"87"),
  2068 => (x"5d",x"5c",x"5b",x"5e"),
  2069 => (x"f4",x"4d",x"71",x"0e"),
  2070 => (x"4a",x"75",x"87",x"e9"),
  2071 => (x"92",x"2a",x"b7",x"c4"),
  2072 => (x"82",x"cc",x"c2",x"c2"),
  2073 => (x"9c",x"cf",x"4c",x"75"),
  2074 => (x"49",x"6a",x"94",x"c2"),
  2075 => (x"c3",x"2b",x"74",x"4b"),
  2076 => (x"74",x"48",x"c2",x"9b"),
  2077 => (x"ff",x"4c",x"70",x"30"),
  2078 => (x"71",x"48",x"74",x"bc"),
  2079 => (x"f3",x"7a",x"70",x"98"),
  2080 => (x"48",x"73",x"87",x"f9"),
  2081 => (x"4c",x"26",x"4d",x"26"),
  2082 => (x"4f",x"26",x"4b",x"26"),
  2083 => (x"00",x"00",x"00",x"00"),
  2084 => (x"00",x"00",x"00",x"00"),
  2085 => (x"00",x"00",x"00",x"00"),
  2086 => (x"00",x"00",x"00",x"00"),
  2087 => (x"00",x"00",x"00",x"00"),
  2088 => (x"00",x"00",x"00",x"00"),
  2089 => (x"00",x"00",x"00",x"00"),
  2090 => (x"00",x"00",x"00",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"00",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"00",x"00"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"00",x"00",x"00",x"00"),
  2096 => (x"00",x"00",x"00",x"00"),
  2097 => (x"00",x"00",x"00",x"00"),
  2098 => (x"00",x"00",x"00",x"00"),
  2099 => (x"48",x"d0",x"ff",x"1e"),
  2100 => (x"71",x"78",x"e1",x"c8"),
  2101 => (x"08",x"d4",x"ff",x"48"),
  2102 => (x"1e",x"4f",x"26",x"78"),
  2103 => (x"c8",x"48",x"d0",x"ff"),
  2104 => (x"48",x"71",x"78",x"e1"),
  2105 => (x"78",x"08",x"d4",x"ff"),
  2106 => (x"ff",x"48",x"66",x"c4"),
  2107 => (x"26",x"78",x"08",x"d4"),
  2108 => (x"4a",x"71",x"1e",x"4f"),
  2109 => (x"1e",x"49",x"66",x"c4"),
  2110 => (x"de",x"ff",x"49",x"72"),
  2111 => (x"48",x"d0",x"ff",x"87"),
  2112 => (x"fc",x"78",x"e0",x"c0"),
  2113 => (x"1e",x"4f",x"26",x"8e"),
  2114 => (x"4b",x"71",x"1e",x"73"),
  2115 => (x"1e",x"49",x"66",x"c8"),
  2116 => (x"e0",x"c1",x"4a",x"73"),
  2117 => (x"d8",x"ff",x"49",x"a2"),
  2118 => (x"26",x"8e",x"fc",x"87"),
  2119 => (x"1e",x"4f",x"26",x"4b"),
  2120 => (x"4b",x"71",x"1e",x"73"),
  2121 => (x"fe",x"49",x"e2",x"c0"),
  2122 => (x"4a",x"c7",x"87",x"e2"),
  2123 => (x"d4",x"ff",x"48",x"13"),
  2124 => (x"49",x"72",x"78",x"08"),
  2125 => (x"99",x"71",x"8a",x"c1"),
  2126 => (x"ff",x"87",x"f1",x"05"),
  2127 => (x"e0",x"c0",x"48",x"d0"),
  2128 => (x"26",x"4b",x"26",x"78"),
  2129 => (x"d0",x"ff",x"1e",x"4f"),
  2130 => (x"78",x"c9",x"c8",x"48"),
  2131 => (x"d4",x"ff",x"48",x"71"),
  2132 => (x"4f",x"26",x"78",x"08"),
  2133 => (x"49",x"4a",x"71",x"1e"),
  2134 => (x"d0",x"ff",x"87",x"eb"),
  2135 => (x"26",x"78",x"c8",x"48"),
  2136 => (x"1e",x"73",x"1e",x"4f"),
  2137 => (x"d1",x"c4",x"4b",x"71"),
  2138 => (x"c3",x"02",x"bf",x"f4"),
  2139 => (x"87",x"eb",x"c2",x"87"),
  2140 => (x"c8",x"48",x"d0",x"ff"),
  2141 => (x"48",x"73",x"78",x"c9"),
  2142 => (x"ff",x"b0",x"e0",x"c0"),
  2143 => (x"c4",x"78",x"08",x"d4"),
  2144 => (x"c0",x"48",x"e8",x"d1"),
  2145 => (x"02",x"66",x"c8",x"78"),
  2146 => (x"ff",x"c3",x"87",x"c5"),
  2147 => (x"c0",x"87",x"c2",x"49"),
  2148 => (x"f0",x"d1",x"c4",x"49"),
  2149 => (x"02",x"66",x"cc",x"59"),
  2150 => (x"d5",x"c5",x"87",x"c6"),
  2151 => (x"87",x"c4",x"4a",x"d5"),
  2152 => (x"4a",x"ff",x"ff",x"cf"),
  2153 => (x"5a",x"f4",x"d1",x"c4"),
  2154 => (x"48",x"f4",x"d1",x"c4"),
  2155 => (x"4b",x"26",x"78",x"c1"),
  2156 => (x"5e",x"0e",x"4f",x"26"),
  2157 => (x"0e",x"5d",x"5c",x"5b"),
  2158 => (x"d1",x"c4",x"4d",x"71"),
  2159 => (x"75",x"4b",x"bf",x"f0"),
  2160 => (x"87",x"cb",x"02",x"9d"),
  2161 => (x"c2",x"91",x"c8",x"49"),
  2162 => (x"71",x"4a",x"d8",x"c5"),
  2163 => (x"c2",x"87",x"c4",x"82"),
  2164 => (x"c0",x"4a",x"d8",x"c9"),
  2165 => (x"73",x"49",x"12",x"4c"),
  2166 => (x"ec",x"d1",x"c4",x"99"),
  2167 => (x"b8",x"71",x"48",x"bf"),
  2168 => (x"78",x"08",x"d4",x"ff"),
  2169 => (x"84",x"2b",x"b7",x"c1"),
  2170 => (x"04",x"ac",x"b7",x"c8"),
  2171 => (x"d1",x"c4",x"87",x"e7"),
  2172 => (x"c8",x"48",x"bf",x"e8"),
  2173 => (x"ec",x"d1",x"c4",x"80"),
  2174 => (x"26",x"4d",x"26",x"58"),
  2175 => (x"26",x"4b",x"26",x"4c"),
  2176 => (x"1e",x"73",x"1e",x"4f"),
  2177 => (x"4a",x"13",x"4b",x"71"),
  2178 => (x"87",x"cb",x"02",x"9a"),
  2179 => (x"e1",x"fe",x"49",x"72"),
  2180 => (x"9a",x"4a",x"13",x"87"),
  2181 => (x"26",x"87",x"f5",x"05"),
  2182 => (x"1e",x"4f",x"26",x"4b"),
  2183 => (x"bf",x"e8",x"d1",x"c4"),
  2184 => (x"e8",x"d1",x"c4",x"49"),
  2185 => (x"78",x"a1",x"c1",x"48"),
  2186 => (x"a9",x"b7",x"c0",x"c4"),
  2187 => (x"ff",x"87",x"db",x"03"),
  2188 => (x"d1",x"c4",x"48",x"d4"),
  2189 => (x"c4",x"78",x"bf",x"ec"),
  2190 => (x"49",x"bf",x"e8",x"d1"),
  2191 => (x"48",x"e8",x"d1",x"c4"),
  2192 => (x"c4",x"78",x"a1",x"c1"),
  2193 => (x"04",x"a9",x"b7",x"c0"),
  2194 => (x"d0",x"ff",x"87",x"e5"),
  2195 => (x"c4",x"78",x"c8",x"48"),
  2196 => (x"c0",x"48",x"f4",x"d1"),
  2197 => (x"00",x"4f",x"26",x"78"),
  2198 => (x"00",x"00",x"00",x"00"),
  2199 => (x"00",x"00",x"00",x"00"),
  2200 => (x"5f",x"00",x"00",x"00"),
  2201 => (x"00",x"00",x"00",x"5f"),
  2202 => (x"00",x"03",x"03",x"00"),
  2203 => (x"00",x"00",x"03",x"03"),
  2204 => (x"14",x"7f",x"7f",x"14"),
  2205 => (x"00",x"14",x"7f",x"7f"),
  2206 => (x"6b",x"2e",x"24",x"00"),
  2207 => (x"00",x"12",x"3a",x"6b"),
  2208 => (x"18",x"36",x"6a",x"4c"),
  2209 => (x"00",x"32",x"56",x"6c"),
  2210 => (x"59",x"4f",x"7e",x"30"),
  2211 => (x"40",x"68",x"3a",x"77"),
  2212 => (x"07",x"04",x"00",x"00"),
  2213 => (x"00",x"00",x"00",x"03"),
  2214 => (x"3e",x"1c",x"00",x"00"),
  2215 => (x"00",x"00",x"41",x"63"),
  2216 => (x"63",x"41",x"00",x"00"),
  2217 => (x"00",x"00",x"1c",x"3e"),
  2218 => (x"1c",x"3e",x"2a",x"08"),
  2219 => (x"08",x"2a",x"3e",x"1c"),
  2220 => (x"3e",x"08",x"08",x"00"),
  2221 => (x"00",x"08",x"08",x"3e"),
  2222 => (x"e0",x"80",x"00",x"00"),
  2223 => (x"00",x"00",x"00",x"60"),
  2224 => (x"08",x"08",x"08",x"00"),
  2225 => (x"00",x"08",x"08",x"08"),
  2226 => (x"60",x"00",x"00",x"00"),
  2227 => (x"00",x"00",x"00",x"60"),
  2228 => (x"18",x"30",x"60",x"40"),
  2229 => (x"01",x"03",x"06",x"0c"),
  2230 => (x"59",x"7f",x"3e",x"00"),
  2231 => (x"00",x"3e",x"7f",x"4d"),
  2232 => (x"7f",x"06",x"04",x"00"),
  2233 => (x"00",x"00",x"00",x"7f"),
  2234 => (x"71",x"63",x"42",x"00"),
  2235 => (x"00",x"46",x"4f",x"59"),
  2236 => (x"49",x"63",x"22",x"00"),
  2237 => (x"00",x"36",x"7f",x"49"),
  2238 => (x"13",x"16",x"1c",x"18"),
  2239 => (x"00",x"10",x"7f",x"7f"),
  2240 => (x"45",x"67",x"27",x"00"),
  2241 => (x"00",x"39",x"7d",x"45"),
  2242 => (x"4b",x"7e",x"3c",x"00"),
  2243 => (x"00",x"30",x"79",x"49"),
  2244 => (x"71",x"01",x"01",x"00"),
  2245 => (x"00",x"07",x"0f",x"79"),
  2246 => (x"49",x"7f",x"36",x"00"),
  2247 => (x"00",x"36",x"7f",x"49"),
  2248 => (x"49",x"4f",x"06",x"00"),
  2249 => (x"00",x"1e",x"3f",x"69"),
  2250 => (x"66",x"00",x"00",x"00"),
  2251 => (x"00",x"00",x"00",x"66"),
  2252 => (x"e6",x"80",x"00",x"00"),
  2253 => (x"00",x"00",x"00",x"66"),
  2254 => (x"14",x"08",x"08",x"00"),
  2255 => (x"00",x"22",x"22",x"14"),
  2256 => (x"14",x"14",x"14",x"00"),
  2257 => (x"00",x"14",x"14",x"14"),
  2258 => (x"14",x"22",x"22",x"00"),
  2259 => (x"00",x"08",x"08",x"14"),
  2260 => (x"51",x"03",x"02",x"00"),
  2261 => (x"00",x"06",x"0f",x"59"),
  2262 => (x"5d",x"41",x"7f",x"3e"),
  2263 => (x"00",x"1e",x"1f",x"55"),
  2264 => (x"09",x"7f",x"7e",x"00"),
  2265 => (x"00",x"7e",x"7f",x"09"),
  2266 => (x"49",x"7f",x"7f",x"00"),
  2267 => (x"00",x"36",x"7f",x"49"),
  2268 => (x"63",x"3e",x"1c",x"00"),
  2269 => (x"00",x"41",x"41",x"41"),
  2270 => (x"41",x"7f",x"7f",x"00"),
  2271 => (x"00",x"1c",x"3e",x"63"),
  2272 => (x"49",x"7f",x"7f",x"00"),
  2273 => (x"00",x"41",x"41",x"49"),
  2274 => (x"09",x"7f",x"7f",x"00"),
  2275 => (x"00",x"01",x"01",x"09"),
  2276 => (x"41",x"7f",x"3e",x"00"),
  2277 => (x"00",x"7a",x"7b",x"49"),
  2278 => (x"08",x"7f",x"7f",x"00"),
  2279 => (x"00",x"7f",x"7f",x"08"),
  2280 => (x"7f",x"41",x"00",x"00"),
  2281 => (x"00",x"00",x"41",x"7f"),
  2282 => (x"40",x"60",x"20",x"00"),
  2283 => (x"00",x"3f",x"7f",x"40"),
  2284 => (x"1c",x"08",x"7f",x"7f"),
  2285 => (x"00",x"41",x"63",x"36"),
  2286 => (x"40",x"7f",x"7f",x"00"),
  2287 => (x"00",x"40",x"40",x"40"),
  2288 => (x"0c",x"06",x"7f",x"7f"),
  2289 => (x"00",x"7f",x"7f",x"06"),
  2290 => (x"0c",x"06",x"7f",x"7f"),
  2291 => (x"00",x"7f",x"7f",x"18"),
  2292 => (x"41",x"7f",x"3e",x"00"),
  2293 => (x"00",x"3e",x"7f",x"41"),
  2294 => (x"09",x"7f",x"7f",x"00"),
  2295 => (x"00",x"06",x"0f",x"09"),
  2296 => (x"61",x"41",x"7f",x"3e"),
  2297 => (x"00",x"40",x"7e",x"7f"),
  2298 => (x"09",x"7f",x"7f",x"00"),
  2299 => (x"00",x"66",x"7f",x"19"),
  2300 => (x"4d",x"6f",x"26",x"00"),
  2301 => (x"00",x"32",x"7b",x"59"),
  2302 => (x"7f",x"01",x"01",x"00"),
  2303 => (x"00",x"01",x"01",x"7f"),
  2304 => (x"40",x"7f",x"3f",x"00"),
  2305 => (x"00",x"3f",x"7f",x"40"),
  2306 => (x"70",x"3f",x"0f",x"00"),
  2307 => (x"00",x"0f",x"3f",x"70"),
  2308 => (x"18",x"30",x"7f",x"7f"),
  2309 => (x"00",x"7f",x"7f",x"30"),
  2310 => (x"1c",x"36",x"63",x"41"),
  2311 => (x"41",x"63",x"36",x"1c"),
  2312 => (x"7c",x"06",x"03",x"01"),
  2313 => (x"01",x"03",x"06",x"7c"),
  2314 => (x"4d",x"59",x"71",x"61"),
  2315 => (x"00",x"41",x"43",x"47"),
  2316 => (x"7f",x"7f",x"00",x"00"),
  2317 => (x"00",x"00",x"41",x"41"),
  2318 => (x"0c",x"06",x"03",x"01"),
  2319 => (x"40",x"60",x"30",x"18"),
  2320 => (x"41",x"41",x"00",x"00"),
  2321 => (x"00",x"00",x"7f",x"7f"),
  2322 => (x"03",x"06",x"0c",x"08"),
  2323 => (x"00",x"08",x"0c",x"06"),
  2324 => (x"80",x"80",x"80",x"80"),
  2325 => (x"00",x"80",x"80",x"80"),
  2326 => (x"03",x"00",x"00",x"00"),
  2327 => (x"00",x"00",x"04",x"07"),
  2328 => (x"54",x"74",x"20",x"00"),
  2329 => (x"00",x"78",x"7c",x"54"),
  2330 => (x"44",x"7f",x"7f",x"00"),
  2331 => (x"00",x"38",x"7c",x"44"),
  2332 => (x"44",x"7c",x"38",x"00"),
  2333 => (x"00",x"00",x"44",x"44"),
  2334 => (x"44",x"7c",x"38",x"00"),
  2335 => (x"00",x"7f",x"7f",x"44"),
  2336 => (x"54",x"7c",x"38",x"00"),
  2337 => (x"00",x"18",x"5c",x"54"),
  2338 => (x"7f",x"7e",x"04",x"00"),
  2339 => (x"00",x"00",x"05",x"05"),
  2340 => (x"a4",x"bc",x"18",x"00"),
  2341 => (x"00",x"7c",x"fc",x"a4"),
  2342 => (x"04",x"7f",x"7f",x"00"),
  2343 => (x"00",x"78",x"7c",x"04"),
  2344 => (x"3d",x"00",x"00",x"00"),
  2345 => (x"00",x"00",x"40",x"7d"),
  2346 => (x"80",x"80",x"80",x"00"),
  2347 => (x"00",x"00",x"7d",x"fd"),
  2348 => (x"10",x"7f",x"7f",x"00"),
  2349 => (x"00",x"44",x"6c",x"38"),
  2350 => (x"3f",x"00",x"00",x"00"),
  2351 => (x"00",x"00",x"40",x"7f"),
  2352 => (x"18",x"0c",x"7c",x"7c"),
  2353 => (x"00",x"78",x"7c",x"0c"),
  2354 => (x"04",x"7c",x"7c",x"00"),
  2355 => (x"00",x"78",x"7c",x"04"),
  2356 => (x"44",x"7c",x"38",x"00"),
  2357 => (x"00",x"38",x"7c",x"44"),
  2358 => (x"24",x"fc",x"fc",x"00"),
  2359 => (x"00",x"18",x"3c",x"24"),
  2360 => (x"24",x"3c",x"18",x"00"),
  2361 => (x"00",x"fc",x"fc",x"24"),
  2362 => (x"04",x"7c",x"7c",x"00"),
  2363 => (x"00",x"08",x"0c",x"04"),
  2364 => (x"54",x"5c",x"48",x"00"),
  2365 => (x"00",x"20",x"74",x"54"),
  2366 => (x"7f",x"3f",x"04",x"00"),
  2367 => (x"00",x"00",x"44",x"44"),
  2368 => (x"40",x"7c",x"3c",x"00"),
  2369 => (x"00",x"7c",x"7c",x"40"),
  2370 => (x"60",x"3c",x"1c",x"00"),
  2371 => (x"00",x"1c",x"3c",x"60"),
  2372 => (x"30",x"60",x"7c",x"3c"),
  2373 => (x"00",x"3c",x"7c",x"60"),
  2374 => (x"10",x"38",x"6c",x"44"),
  2375 => (x"00",x"44",x"6c",x"38"),
  2376 => (x"e0",x"bc",x"1c",x"00"),
  2377 => (x"00",x"1c",x"3c",x"60"),
  2378 => (x"74",x"64",x"44",x"00"),
  2379 => (x"00",x"44",x"4c",x"5c"),
  2380 => (x"3e",x"08",x"08",x"00"),
  2381 => (x"00",x"41",x"41",x"77"),
  2382 => (x"7f",x"00",x"00",x"00"),
  2383 => (x"00",x"00",x"00",x"7f"),
  2384 => (x"77",x"41",x"41",x"00"),
  2385 => (x"00",x"08",x"08",x"3e"),
  2386 => (x"03",x"01",x"01",x"02"),
  2387 => (x"00",x"01",x"02",x"02"),
  2388 => (x"7f",x"7f",x"7f",x"7f"),
  2389 => (x"00",x"7f",x"7f",x"7f"),
  2390 => (x"1c",x"1c",x"08",x"08"),
  2391 => (x"7f",x"7f",x"3e",x"3e"),
  2392 => (x"3e",x"3e",x"7f",x"7f"),
  2393 => (x"08",x"08",x"1c",x"1c"),
  2394 => (x"7c",x"18",x"10",x"00"),
  2395 => (x"00",x"10",x"18",x"7c"),
  2396 => (x"7c",x"30",x"10",x"00"),
  2397 => (x"00",x"10",x"30",x"7c"),
  2398 => (x"60",x"60",x"30",x"10"),
  2399 => (x"00",x"06",x"1e",x"78"),
  2400 => (x"18",x"3c",x"66",x"42"),
  2401 => (x"00",x"42",x"66",x"3c"),
  2402 => (x"c2",x"6a",x"38",x"78"),
  2403 => (x"00",x"38",x"6c",x"c6"),
  2404 => (x"60",x"00",x"00",x"60"),
  2405 => (x"00",x"60",x"00",x"00"),
  2406 => (x"5c",x"5b",x"5e",x"0e"),
  2407 => (x"86",x"fc",x"0e",x"5d"),
  2408 => (x"d2",x"c4",x"7e",x"71"),
  2409 => (x"c0",x"4c",x"bf",x"c8"),
  2410 => (x"c4",x"1e",x"c0",x"4b"),
  2411 => (x"c4",x"02",x"ab",x"66"),
  2412 => (x"c2",x"4d",x"c0",x"87"),
  2413 => (x"75",x"4d",x"c1",x"87"),
  2414 => (x"ee",x"49",x"73",x"1e"),
  2415 => (x"86",x"c8",x"87",x"e3"),
  2416 => (x"ef",x"49",x"e0",x"c0"),
  2417 => (x"a4",x"c4",x"87",x"ec"),
  2418 => (x"f0",x"49",x"6a",x"4a"),
  2419 => (x"ca",x"f1",x"87",x"f3"),
  2420 => (x"c1",x"84",x"cc",x"87"),
  2421 => (x"ab",x"b7",x"c8",x"83"),
  2422 => (x"87",x"cd",x"ff",x"04"),
  2423 => (x"4d",x"26",x"8e",x"fc"),
  2424 => (x"4b",x"26",x"4c",x"26"),
  2425 => (x"71",x"1e",x"4f",x"26"),
  2426 => (x"cc",x"d2",x"c4",x"4a"),
  2427 => (x"cc",x"d2",x"c4",x"5a"),
  2428 => (x"49",x"78",x"c7",x"48"),
  2429 => (x"26",x"87",x"e1",x"fe"),
  2430 => (x"1e",x"73",x"1e",x"4f"),
  2431 => (x"b7",x"c0",x"4a",x"71"),
  2432 => (x"87",x"d3",x"03",x"aa"),
  2433 => (x"bf",x"d4",x"e6",x"c2"),
  2434 => (x"c1",x"87",x"c4",x"05"),
  2435 => (x"c0",x"87",x"c2",x"4b"),
  2436 => (x"d8",x"e6",x"c2",x"4b"),
  2437 => (x"c2",x"87",x"c4",x"5b"),
  2438 => (x"c2",x"5a",x"d8",x"e6"),
  2439 => (x"4a",x"bf",x"d4",x"e6"),
  2440 => (x"c0",x"c1",x"9a",x"c1"),
  2441 => (x"eb",x"ec",x"49",x"a2"),
  2442 => (x"c2",x"48",x"fc",x"87"),
  2443 => (x"78",x"bf",x"d4",x"e6"),
  2444 => (x"4f",x"26",x"4b",x"26"),
  2445 => (x"d4",x"e6",x"c2",x"1e"),
  2446 => (x"4f",x"26",x"48",x"bf"),
  2447 => (x"c4",x"4a",x"71",x"1e"),
  2448 => (x"49",x"72",x"1e",x"66"),
  2449 => (x"fc",x"87",x"c0",x"eb"),
  2450 => (x"1e",x"4f",x"26",x"8e"),
  2451 => (x"c3",x"48",x"d4",x"ff"),
  2452 => (x"d0",x"ff",x"78",x"ff"),
  2453 => (x"78",x"e1",x"c0",x"48"),
  2454 => (x"c1",x"48",x"d4",x"ff"),
  2455 => (x"c4",x"48",x"71",x"78"),
  2456 => (x"08",x"d4",x"ff",x"30"),
  2457 => (x"48",x"d0",x"ff",x"78"),
  2458 => (x"26",x"78",x"e0",x"c0"),
  2459 => (x"e6",x"c2",x"1e",x"4f"),
  2460 => (x"c1",x"49",x"bf",x"d4"),
  2461 => (x"c4",x"87",x"f5",x"d4"),
  2462 => (x"e8",x"48",x"c0",x"d2"),
  2463 => (x"d1",x"c4",x"78",x"bf"),
  2464 => (x"bf",x"ec",x"48",x"fc"),
  2465 => (x"c0",x"d2",x"c4",x"78"),
  2466 => (x"c3",x"49",x"4a",x"bf"),
  2467 => (x"b7",x"c8",x"99",x"ff"),
  2468 => (x"71",x"48",x"72",x"2a"),
  2469 => (x"c8",x"d2",x"c4",x"b0"),
  2470 => (x"0e",x"4f",x"26",x"58"),
  2471 => (x"5d",x"5c",x"5b",x"5e"),
  2472 => (x"ff",x"4b",x"71",x"0e"),
  2473 => (x"d1",x"c4",x"87",x"c7"),
  2474 => (x"50",x"c0",x"48",x"f8"),
  2475 => (x"de",x"e6",x"49",x"73"),
  2476 => (x"4c",x"49",x"70",x"87"),
  2477 => (x"ee",x"cb",x"9c",x"c2"),
  2478 => (x"87",x"e0",x"cb",x"49"),
  2479 => (x"d1",x"c4",x"4d",x"70"),
  2480 => (x"05",x"bf",x"97",x"f8"),
  2481 => (x"d0",x"87",x"e2",x"c1"),
  2482 => (x"d2",x"c4",x"49",x"66"),
  2483 => (x"05",x"99",x"bf",x"c4"),
  2484 => (x"66",x"d4",x"87",x"d6"),
  2485 => (x"fc",x"d1",x"c4",x"49"),
  2486 => (x"cb",x"05",x"99",x"bf"),
  2487 => (x"e5",x"49",x"73",x"87"),
  2488 => (x"98",x"70",x"87",x"ed"),
  2489 => (x"87",x"c1",x"c1",x"02"),
  2490 => (x"c0",x"fe",x"4c",x"c1"),
  2491 => (x"ca",x"49",x"75",x"87"),
  2492 => (x"98",x"70",x"87",x"f6"),
  2493 => (x"c4",x"87",x"c6",x"02"),
  2494 => (x"c1",x"48",x"f8",x"d1"),
  2495 => (x"f8",x"d1",x"c4",x"50"),
  2496 => (x"c0",x"05",x"bf",x"97"),
  2497 => (x"d2",x"c4",x"87",x"e3"),
  2498 => (x"d0",x"49",x"bf",x"c4"),
  2499 => (x"ff",x"05",x"99",x"66"),
  2500 => (x"d1",x"c4",x"87",x"d6"),
  2501 => (x"d4",x"49",x"bf",x"fc"),
  2502 => (x"ff",x"05",x"99",x"66"),
  2503 => (x"49",x"73",x"87",x"ca"),
  2504 => (x"70",x"87",x"ec",x"e4"),
  2505 => (x"ff",x"fe",x"05",x"98"),
  2506 => (x"26",x"48",x"74",x"87"),
  2507 => (x"26",x"4c",x"26",x"4d"),
  2508 => (x"0e",x"4f",x"26",x"4b"),
  2509 => (x"5d",x"5c",x"5b",x"5e"),
  2510 => (x"c0",x"86",x"f8",x"0e"),
  2511 => (x"bf",x"ec",x"4c",x"4d"),
  2512 => (x"48",x"a6",x"c4",x"7e"),
  2513 => (x"bf",x"c8",x"d2",x"c4"),
  2514 => (x"c0",x"1e",x"c1",x"78"),
  2515 => (x"fd",x"49",x"c7",x"1e"),
  2516 => (x"86",x"c8",x"87",x"c9"),
  2517 => (x"cd",x"02",x"98",x"70"),
  2518 => (x"fa",x"49",x"ff",x"87"),
  2519 => (x"da",x"c1",x"87",x"db"),
  2520 => (x"87",x"eb",x"e3",x"49"),
  2521 => (x"d1",x"c4",x"4d",x"c1"),
  2522 => (x"02",x"bf",x"97",x"f8"),
  2523 => (x"e6",x"c2",x"87",x"cf"),
  2524 => (x"c1",x"49",x"bf",x"cc"),
  2525 => (x"d0",x"e6",x"c2",x"b9"),
  2526 => (x"ce",x"fb",x"71",x"59"),
  2527 => (x"c0",x"d2",x"c4",x"87"),
  2528 => (x"e6",x"c2",x"4b",x"bf"),
  2529 => (x"c0",x"05",x"bf",x"d4"),
  2530 => (x"fd",x"c3",x"87",x"e9"),
  2531 => (x"87",x"ff",x"e2",x"49"),
  2532 => (x"e2",x"49",x"fa",x"c3"),
  2533 => (x"49",x"73",x"87",x"f9"),
  2534 => (x"71",x"99",x"ff",x"c3"),
  2535 => (x"fa",x"49",x"c0",x"1e"),
  2536 => (x"49",x"73",x"87",x"da"),
  2537 => (x"71",x"29",x"b7",x"c8"),
  2538 => (x"fa",x"49",x"c1",x"1e"),
  2539 => (x"86",x"c8",x"87",x"ce"),
  2540 => (x"c4",x"87",x"f4",x"c5"),
  2541 => (x"4b",x"bf",x"c4",x"d2"),
  2542 => (x"87",x"dd",x"02",x"9b"),
  2543 => (x"bf",x"d0",x"e6",x"c2"),
  2544 => (x"87",x"e4",x"c7",x"49"),
  2545 => (x"c4",x"05",x"98",x"70"),
  2546 => (x"d2",x"4b",x"c0",x"87"),
  2547 => (x"49",x"e0",x"c2",x"87"),
  2548 => (x"c2",x"87",x"c9",x"c7"),
  2549 => (x"c6",x"58",x"d4",x"e6"),
  2550 => (x"d0",x"e6",x"c2",x"87"),
  2551 => (x"73",x"78",x"c0",x"48"),
  2552 => (x"05",x"99",x"c2",x"49"),
  2553 => (x"eb",x"c3",x"87",x"cd"),
  2554 => (x"87",x"e3",x"e1",x"49"),
  2555 => (x"99",x"c2",x"49",x"70"),
  2556 => (x"fb",x"87",x"c2",x"02"),
  2557 => (x"c1",x"49",x"73",x"4c"),
  2558 => (x"87",x"cd",x"05",x"99"),
  2559 => (x"e1",x"49",x"f4",x"c3"),
  2560 => (x"49",x"70",x"87",x"cd"),
  2561 => (x"c2",x"02",x"99",x"c2"),
  2562 => (x"73",x"4c",x"fa",x"87"),
  2563 => (x"05",x"99",x"c8",x"49"),
  2564 => (x"f5",x"c3",x"87",x"cd"),
  2565 => (x"87",x"f7",x"e0",x"49"),
  2566 => (x"99",x"c2",x"49",x"70"),
  2567 => (x"c4",x"87",x"d5",x"02"),
  2568 => (x"02",x"bf",x"cc",x"d2"),
  2569 => (x"c1",x"48",x"87",x"ca"),
  2570 => (x"d0",x"d2",x"c4",x"88"),
  2571 => (x"87",x"c2",x"c0",x"58"),
  2572 => (x"4d",x"c1",x"4c",x"ff"),
  2573 => (x"99",x"c4",x"49",x"73"),
  2574 => (x"c3",x"87",x"cd",x"05"),
  2575 => (x"ce",x"e0",x"49",x"f2"),
  2576 => (x"c2",x"49",x"70",x"87"),
  2577 => (x"87",x"dc",x"02",x"99"),
  2578 => (x"bf",x"cc",x"d2",x"c4"),
  2579 => (x"b7",x"c7",x"48",x"7e"),
  2580 => (x"cb",x"c0",x"03",x"a8"),
  2581 => (x"c1",x"48",x"6e",x"87"),
  2582 => (x"d0",x"d2",x"c4",x"80"),
  2583 => (x"87",x"c2",x"c0",x"58"),
  2584 => (x"4d",x"c1",x"4c",x"fe"),
  2585 => (x"ff",x"49",x"fd",x"c3"),
  2586 => (x"70",x"87",x"e4",x"df"),
  2587 => (x"02",x"99",x"c2",x"49"),
  2588 => (x"d2",x"c4",x"87",x"d5"),
  2589 => (x"c0",x"02",x"bf",x"cc"),
  2590 => (x"d2",x"c4",x"87",x"c9"),
  2591 => (x"78",x"c0",x"48",x"cc"),
  2592 => (x"fd",x"87",x"c2",x"c0"),
  2593 => (x"c3",x"4d",x"c1",x"4c"),
  2594 => (x"df",x"ff",x"49",x"fa"),
  2595 => (x"49",x"70",x"87",x"c1"),
  2596 => (x"c0",x"02",x"99",x"c2"),
  2597 => (x"d2",x"c4",x"87",x"d9"),
  2598 => (x"c7",x"48",x"bf",x"cc"),
  2599 => (x"c0",x"03",x"a8",x"b7"),
  2600 => (x"d2",x"c4",x"87",x"c9"),
  2601 => (x"78",x"c7",x"48",x"cc"),
  2602 => (x"fc",x"87",x"c2",x"c0"),
  2603 => (x"c0",x"4d",x"c1",x"4c"),
  2604 => (x"c0",x"03",x"ac",x"b7"),
  2605 => (x"66",x"c4",x"87",x"d3"),
  2606 => (x"80",x"e0",x"c1",x"48"),
  2607 => (x"bf",x"6e",x"7e",x"70"),
  2608 => (x"87",x"c5",x"c0",x"02"),
  2609 => (x"73",x"49",x"74",x"4b"),
  2610 => (x"c3",x"1e",x"c0",x"0f"),
  2611 => (x"da",x"c1",x"1e",x"f0"),
  2612 => (x"87",x"c7",x"f7",x"49"),
  2613 => (x"98",x"70",x"86",x"c8"),
  2614 => (x"87",x"d8",x"c0",x"02"),
  2615 => (x"bf",x"cc",x"d2",x"c4"),
  2616 => (x"cc",x"49",x"6e",x"7e"),
  2617 => (x"4a",x"66",x"c4",x"91"),
  2618 => (x"02",x"6a",x"82",x"71"),
  2619 => (x"4b",x"87",x"c5",x"c0"),
  2620 => (x"0f",x"73",x"49",x"6e"),
  2621 => (x"c0",x"02",x"9d",x"75"),
  2622 => (x"d2",x"c4",x"87",x"c8"),
  2623 => (x"f2",x"49",x"bf",x"cc"),
  2624 => (x"e6",x"c2",x"87",x"d6"),
  2625 => (x"c0",x"02",x"bf",x"d8"),
  2626 => (x"c2",x"49",x"87",x"dd"),
  2627 => (x"98",x"70",x"87",x"da"),
  2628 => (x"87",x"d3",x"c0",x"02"),
  2629 => (x"bf",x"cc",x"d2",x"c4"),
  2630 => (x"87",x"fc",x"f1",x"49"),
  2631 => (x"d8",x"f3",x"49",x"c0"),
  2632 => (x"d8",x"e6",x"c2",x"87"),
  2633 => (x"f8",x"78",x"c0",x"48"),
  2634 => (x"26",x"4d",x"26",x"8e"),
  2635 => (x"26",x"4b",x"26",x"4c"),
  2636 => (x"5b",x"5e",x"0e",x"4f"),
  2637 => (x"fc",x"0e",x"5d",x"5c"),
  2638 => (x"c4",x"4c",x"71",x"86"),
  2639 => (x"49",x"bf",x"c8",x"d2"),
  2640 => (x"4d",x"a1",x"d4",x"c1"),
  2641 => (x"69",x"81",x"d8",x"c1"),
  2642 => (x"02",x"9c",x"74",x"7e"),
  2643 => (x"a5",x"c4",x"87",x"cf"),
  2644 => (x"c4",x"7b",x"74",x"4b"),
  2645 => (x"49",x"bf",x"c8",x"d2"),
  2646 => (x"6e",x"87",x"cb",x"f2"),
  2647 => (x"05",x"9c",x"74",x"7b"),
  2648 => (x"4b",x"c0",x"87",x"c4"),
  2649 => (x"4b",x"c1",x"87",x"c2"),
  2650 => (x"cc",x"f2",x"49",x"73"),
  2651 => (x"02",x"66",x"d4",x"87"),
  2652 => (x"c0",x"49",x"87",x"c8"),
  2653 => (x"4a",x"70",x"87",x"e6"),
  2654 => (x"4a",x"c0",x"87",x"c2"),
  2655 => (x"5a",x"dc",x"e6",x"c2"),
  2656 => (x"4d",x"26",x"8e",x"fc"),
  2657 => (x"4b",x"26",x"4c",x"26"),
  2658 => (x"00",x"00",x"4f",x"26"),
  2659 => (x"00",x"00",x"00",x"00"),
  2660 => (x"00",x"00",x"00",x"00"),
  2661 => (x"00",x"00",x"00",x"00"),
  2662 => (x"00",x"00",x"00",x"00"),
  2663 => (x"ff",x"4a",x"71",x"1e"),
  2664 => (x"72",x"49",x"bf",x"c8"),
  2665 => (x"4f",x"26",x"48",x"a1"),
  2666 => (x"bf",x"c8",x"ff",x"1e"),
  2667 => (x"c0",x"c0",x"fe",x"89"),
  2668 => (x"a9",x"c0",x"c0",x"c0"),
  2669 => (x"c0",x"87",x"c4",x"01"),
  2670 => (x"c1",x"87",x"c2",x"4a"),
  2671 => (x"26",x"48",x"72",x"4a"),
  2672 => (x"5b",x"5e",x"0e",x"4f"),
  2673 => (x"71",x"0e",x"5d",x"5c"),
  2674 => (x"4c",x"d4",x"ff",x"4b"),
  2675 => (x"c0",x"48",x"66",x"d0"),
  2676 => (x"ff",x"49",x"d6",x"78"),
  2677 => (x"c3",x"87",x"f5",x"db"),
  2678 => (x"49",x"6c",x"7c",x"ff"),
  2679 => (x"71",x"99",x"ff",x"c3"),
  2680 => (x"f0",x"c3",x"49",x"4d"),
  2681 => (x"a9",x"e0",x"c1",x"99"),
  2682 => (x"c3",x"87",x"cb",x"05"),
  2683 => (x"48",x"6c",x"7c",x"ff"),
  2684 => (x"66",x"d0",x"98",x"c3"),
  2685 => (x"ff",x"c3",x"78",x"08"),
  2686 => (x"49",x"4a",x"6c",x"7c"),
  2687 => (x"ff",x"c3",x"31",x"c8"),
  2688 => (x"71",x"4a",x"6c",x"7c"),
  2689 => (x"c8",x"49",x"72",x"b2"),
  2690 => (x"7c",x"ff",x"c3",x"31"),
  2691 => (x"b2",x"71",x"4a",x"6c"),
  2692 => (x"31",x"c8",x"49",x"72"),
  2693 => (x"6c",x"7c",x"ff",x"c3"),
  2694 => (x"ff",x"b2",x"71",x"4a"),
  2695 => (x"e0",x"c0",x"48",x"d0"),
  2696 => (x"02",x"9b",x"73",x"78"),
  2697 => (x"7b",x"72",x"87",x"c2"),
  2698 => (x"4d",x"26",x"48",x"75"),
  2699 => (x"4b",x"26",x"4c",x"26"),
  2700 => (x"26",x"1e",x"4f",x"26"),
  2701 => (x"5b",x"5e",x"0e",x"4f"),
  2702 => (x"86",x"f8",x"0e",x"5c"),
  2703 => (x"a6",x"c8",x"1e",x"76"),
  2704 => (x"87",x"fd",x"fd",x"49"),
  2705 => (x"4b",x"70",x"86",x"c4"),
  2706 => (x"a8",x"c4",x"48",x"6e"),
  2707 => (x"87",x"f4",x"c2",x"03"),
  2708 => (x"f0",x"c3",x"4a",x"73"),
  2709 => (x"aa",x"d0",x"c1",x"9a"),
  2710 => (x"c1",x"87",x"c7",x"02"),
  2711 => (x"c2",x"05",x"aa",x"e0"),
  2712 => (x"49",x"73",x"87",x"e2"),
  2713 => (x"c3",x"02",x"99",x"c8"),
  2714 => (x"87",x"c6",x"ff",x"87"),
  2715 => (x"9c",x"c3",x"4c",x"73"),
  2716 => (x"c1",x"05",x"ac",x"c2"),
  2717 => (x"66",x"c4",x"87",x"c4"),
  2718 => (x"71",x"31",x"c9",x"49"),
  2719 => (x"4a",x"66",x"c4",x"1e"),
  2720 => (x"c4",x"92",x"c8",x"c1"),
  2721 => (x"72",x"49",x"d0",x"d2"),
  2722 => (x"fe",x"c3",x"fe",x"81"),
  2723 => (x"ff",x"49",x"d8",x"87"),
  2724 => (x"c8",x"87",x"f9",x"d8"),
  2725 => (x"ff",x"c3",x"1e",x"c0"),
  2726 => (x"db",x"fd",x"49",x"d0"),
  2727 => (x"d0",x"ff",x"87",x"c9"),
  2728 => (x"78",x"e0",x"c0",x"48"),
  2729 => (x"1e",x"d0",x"ff",x"c3"),
  2730 => (x"c1",x"4a",x"66",x"cc"),
  2731 => (x"d2",x"c4",x"92",x"c8"),
  2732 => (x"81",x"72",x"49",x"d0"),
  2733 => (x"87",x"c8",x"ff",x"fd"),
  2734 => (x"ac",x"c1",x"86",x"cc"),
  2735 => (x"87",x"c4",x"c1",x"05"),
  2736 => (x"c9",x"49",x"66",x"c4"),
  2737 => (x"c4",x"1e",x"71",x"31"),
  2738 => (x"c8",x"c1",x"4a",x"66"),
  2739 => (x"d0",x"d2",x"c4",x"92"),
  2740 => (x"fe",x"81",x"72",x"49"),
  2741 => (x"c3",x"87",x"f4",x"c2"),
  2742 => (x"c8",x"1e",x"d0",x"ff"),
  2743 => (x"c8",x"c1",x"4a",x"66"),
  2744 => (x"d0",x"d2",x"c4",x"92"),
  2745 => (x"fd",x"81",x"72",x"49"),
  2746 => (x"d7",x"87",x"c6",x"fd"),
  2747 => (x"db",x"d7",x"ff",x"49"),
  2748 => (x"1e",x"c0",x"c8",x"87"),
  2749 => (x"49",x"d0",x"ff",x"c3"),
  2750 => (x"87",x"c8",x"d9",x"fd"),
  2751 => (x"d0",x"ff",x"86",x"cc"),
  2752 => (x"78",x"e0",x"c0",x"48"),
  2753 => (x"4c",x"26",x"8e",x"f8"),
  2754 => (x"4f",x"26",x"4b",x"26"),
  2755 => (x"5c",x"5b",x"5e",x"0e"),
  2756 => (x"4a",x"71",x"0e",x"5d"),
  2757 => (x"d0",x"4c",x"d4",x"ff"),
  2758 => (x"b7",x"c3",x"4d",x"66"),
  2759 => (x"87",x"c5",x"06",x"ad"),
  2760 => (x"e2",x"c1",x"48",x"c0"),
  2761 => (x"75",x"1e",x"72",x"87"),
  2762 => (x"93",x"c8",x"c1",x"4b"),
  2763 => (x"83",x"d0",x"d2",x"c4"),
  2764 => (x"f5",x"fd",x"49",x"73"),
  2765 => (x"83",x"c8",x"87",x"fd"),
  2766 => (x"d0",x"ff",x"4b",x"6b"),
  2767 => (x"78",x"e1",x"c8",x"48"),
  2768 => (x"48",x"73",x"7c",x"dd"),
  2769 => (x"70",x"98",x"ff",x"c3"),
  2770 => (x"c8",x"49",x"73",x"7c"),
  2771 => (x"48",x"71",x"29",x"b7"),
  2772 => (x"70",x"98",x"ff",x"c3"),
  2773 => (x"d0",x"49",x"73",x"7c"),
  2774 => (x"48",x"71",x"29",x"b7"),
  2775 => (x"70",x"98",x"ff",x"c3"),
  2776 => (x"d8",x"48",x"73",x"7c"),
  2777 => (x"7c",x"70",x"28",x"b7"),
  2778 => (x"7c",x"7c",x"7c",x"c0"),
  2779 => (x"7c",x"7c",x"7c",x"7c"),
  2780 => (x"7c",x"7c",x"7c",x"7c"),
  2781 => (x"48",x"d0",x"ff",x"7c"),
  2782 => (x"75",x"78",x"e0",x"c0"),
  2783 => (x"ff",x"49",x"dc",x"1e"),
  2784 => (x"c8",x"87",x"ee",x"d5"),
  2785 => (x"26",x"48",x"73",x"86"),
  2786 => (x"26",x"4c",x"26",x"4d"),
  2787 => (x"1e",x"4f",x"26",x"4b"),
  2788 => (x"86",x"fc",x"1e",x"73"),
  2789 => (x"f0",x"c0",x"4b",x"71"),
  2790 => (x"ec",x"c0",x"4a",x"a3"),
  2791 => (x"82",x"69",x"49",x"a3"),
  2792 => (x"69",x"52",x"66",x"cc"),
  2793 => (x"70",x"80",x"c1",x"48"),
  2794 => (x"98",x"cf",x"48",x"7e"),
  2795 => (x"8e",x"fc",x"79",x"70"),
  2796 => (x"4f",x"26",x"4b",x"26"),
  2797 => (x"5c",x"5b",x"5e",x"0e"),
  2798 => (x"e9",x"4b",x"71",x"0e"),
  2799 => (x"4c",x"70",x"87",x"f6"),
  2800 => (x"87",x"ff",x"c6",x"ff"),
  2801 => (x"c2",x"49",x"66",x"cc"),
  2802 => (x"dc",x"02",x"99",x"c0"),
  2803 => (x"05",x"9c",x"74",x"87"),
  2804 => (x"e0",x"c3",x"87",x"ca"),
  2805 => (x"fe",x"49",x"73",x"1e"),
  2806 => (x"86",x"c4",x"87",x"f5"),
  2807 => (x"c4",x"1e",x"e0",x"c3"),
  2808 => (x"ff",x"49",x"fc",x"d0"),
  2809 => (x"c4",x"87",x"c2",x"ca"),
  2810 => (x"49",x"66",x"cc",x"86"),
  2811 => (x"02",x"99",x"c0",x"c4"),
  2812 => (x"9c",x"74",x"87",x"dc"),
  2813 => (x"c3",x"87",x"ca",x"05"),
  2814 => (x"49",x"73",x"1e",x"f0"),
  2815 => (x"c4",x"87",x"d0",x"fe"),
  2816 => (x"1e",x"f0",x"c3",x"86"),
  2817 => (x"49",x"fc",x"d0",x"c4"),
  2818 => (x"87",x"dd",x"c9",x"ff"),
  2819 => (x"9c",x"74",x"86",x"c4"),
  2820 => (x"cc",x"87",x"cf",x"05"),
  2821 => (x"ff",x"c1",x"49",x"66"),
  2822 => (x"73",x"1e",x"71",x"99"),
  2823 => (x"87",x"ef",x"fd",x"49"),
  2824 => (x"66",x"cc",x"86",x"c4"),
  2825 => (x"99",x"ff",x"c1",x"49"),
  2826 => (x"d0",x"c4",x"1e",x"71"),
  2827 => (x"c8",x"ff",x"49",x"fc"),
  2828 => (x"c5",x"ff",x"87",x"f7"),
  2829 => (x"8e",x"fc",x"87",x"c5"),
  2830 => (x"4b",x"26",x"4c",x"26"),
  2831 => (x"5e",x"0e",x"4f",x"26"),
  2832 => (x"fc",x"0e",x"5c",x"5b"),
  2833 => (x"fa",x"c4",x"ff",x"86"),
  2834 => (x"c0",x"f3",x"c2",x"87"),
  2835 => (x"d7",x"f5",x"49",x"bf"),
  2836 => (x"02",x"98",x"70",x"87"),
  2837 => (x"c4",x"87",x"dc",x"c1"),
  2838 => (x"48",x"bf",x"dc",x"d7"),
  2839 => (x"bf",x"e0",x"d7",x"c4"),
  2840 => (x"ce",x"c1",x"02",x"a8"),
  2841 => (x"e4",x"d7",x"c4",x"87"),
  2842 => (x"dc",x"d7",x"c4",x"49"),
  2843 => (x"4c",x"11",x"81",x"bf"),
  2844 => (x"aa",x"e0",x"c3",x"4a"),
  2845 => (x"c3",x"87",x"c6",x"02"),
  2846 => (x"c4",x"05",x"aa",x"f0"),
  2847 => (x"c2",x"4b",x"c4",x"87"),
  2848 => (x"73",x"4b",x"cf",x"87"),
  2849 => (x"87",x"d4",x"f4",x"49"),
  2850 => (x"58",x"c4",x"f3",x"c2"),
  2851 => (x"c8",x"48",x"d0",x"ff"),
  2852 => (x"d4",x"ff",x"78",x"e1"),
  2853 => (x"74",x"78",x"c5",x"48"),
  2854 => (x"08",x"d4",x"ff",x"48"),
  2855 => (x"48",x"d0",x"ff",x"78"),
  2856 => (x"c4",x"78",x"e0",x"c0"),
  2857 => (x"48",x"bf",x"dc",x"d7"),
  2858 => (x"7e",x"70",x"80",x"c1"),
  2859 => (x"c4",x"98",x"cf",x"48"),
  2860 => (x"ff",x"58",x"e0",x"d7"),
  2861 => (x"fc",x"87",x"c4",x"c3"),
  2862 => (x"26",x"4c",x"26",x"8e"),
  2863 => (x"00",x"4f",x"26",x"4b"),
  2864 => (x"00",x"00",x"00",x"00"),
  2865 => (x"5c",x"5b",x"5e",x"0e"),
  2866 => (x"dc",x"ff",x"0e",x"5d"),
  2867 => (x"c4",x"7e",x"c0",x"86"),
  2868 => (x"49",x"bf",x"f8",x"d6"),
  2869 => (x"1e",x"71",x"81",x"c2"),
  2870 => (x"4a",x"c6",x"1e",x"72"),
  2871 => (x"87",x"f3",x"d0",x"fd"),
  2872 => (x"4a",x"26",x"48",x"71"),
  2873 => (x"a6",x"cc",x"49",x"26"),
  2874 => (x"f8",x"d6",x"c4",x"58"),
  2875 => (x"81",x"c4",x"49",x"bf"),
  2876 => (x"1e",x"72",x"1e",x"71"),
  2877 => (x"d0",x"fd",x"4a",x"c6"),
  2878 => (x"48",x"71",x"87",x"d9"),
  2879 => (x"49",x"26",x"4a",x"26"),
  2880 => (x"fc",x"58",x"a6",x"d0"),
  2881 => (x"fe",x"c2",x"87",x"f8"),
  2882 => (x"f2",x"49",x"bf",x"d4"),
  2883 => (x"98",x"70",x"87",x"da"),
  2884 => (x"87",x"f4",x"c9",x"02"),
  2885 => (x"f2",x"49",x"e0",x"c0"),
  2886 => (x"fe",x"c2",x"87",x"c2"),
  2887 => (x"4c",x"c0",x"58",x"d8"),
  2888 => (x"91",x"c4",x"49",x"74"),
  2889 => (x"69",x"81",x"d0",x"fe"),
  2890 => (x"c4",x"49",x"74",x"4a"),
  2891 => (x"81",x"bf",x"f8",x"d6"),
  2892 => (x"d7",x"c4",x"91",x"c4"),
  2893 => (x"79",x"72",x"81",x"c4"),
  2894 => (x"87",x"d2",x"02",x"9a"),
  2895 => (x"89",x"c1",x"49",x"72"),
  2896 => (x"48",x"6e",x"9a",x"71"),
  2897 => (x"7e",x"70",x"80",x"c1"),
  2898 => (x"ff",x"05",x"9a",x"72"),
  2899 => (x"84",x"c1",x"87",x"ee"),
  2900 => (x"04",x"ac",x"b7",x"c2"),
  2901 => (x"6e",x"87",x"c9",x"ff"),
  2902 => (x"b7",x"fc",x"c0",x"48"),
  2903 => (x"e7",x"c8",x"04",x"a8"),
  2904 => (x"74",x"4c",x"c0",x"87"),
  2905 => (x"82",x"66",x"c8",x"4a"),
  2906 => (x"d7",x"c4",x"92",x"c4"),
  2907 => (x"49",x"74",x"82",x"c4"),
  2908 => (x"c4",x"81",x"66",x"cc"),
  2909 => (x"c4",x"d7",x"c4",x"91"),
  2910 => (x"69",x"4a",x"6a",x"81"),
  2911 => (x"74",x"b9",x"72",x"49"),
  2912 => (x"f8",x"d6",x"c4",x"4b"),
  2913 => (x"93",x"c4",x"83",x"bf"),
  2914 => (x"83",x"c4",x"d7",x"c4"),
  2915 => (x"48",x"72",x"ba",x"6b"),
  2916 => (x"a6",x"d8",x"98",x"71"),
  2917 => (x"c4",x"49",x"74",x"58"),
  2918 => (x"81",x"bf",x"f8",x"d6"),
  2919 => (x"d7",x"c4",x"91",x"c4"),
  2920 => (x"7e",x"69",x"81",x"c4"),
  2921 => (x"c0",x"48",x"a6",x"d8"),
  2922 => (x"5c",x"a6",x"d4",x"78"),
  2923 => (x"df",x"49",x"66",x"d4"),
  2924 => (x"e2",x"c6",x"02",x"29"),
  2925 => (x"4a",x"66",x"d0",x"87"),
  2926 => (x"d8",x"92",x"e0",x"c0"),
  2927 => (x"ff",x"c0",x"82",x"66"),
  2928 => (x"70",x"88",x"72",x"48"),
  2929 => (x"48",x"a6",x"dc",x"4a"),
  2930 => (x"80",x"c4",x"78",x"c0"),
  2931 => (x"49",x"6e",x"78",x"c0"),
  2932 => (x"4c",x"71",x"29",x"df"),
  2933 => (x"48",x"f4",x"d6",x"c4"),
  2934 => (x"49",x"72",x"78",x"c1"),
  2935 => (x"2a",x"b7",x"31",x"c3"),
  2936 => (x"ff",x"c0",x"b1",x"72"),
  2937 => (x"c3",x"91",x"c4",x"99"),
  2938 => (x"71",x"4d",x"c8",x"f0"),
  2939 => (x"49",x"4b",x"6d",x"85"),
  2940 => (x"99",x"c0",x"c0",x"c4"),
  2941 => (x"74",x"87",x"d6",x"02"),
  2942 => (x"c7",x"c0",x"02",x"9c"),
  2943 => (x"c0",x"80",x"c8",x"87"),
  2944 => (x"87",x"d3",x"c5",x"78"),
  2945 => (x"48",x"fc",x"d6",x"c4"),
  2946 => (x"ca",x"c5",x"78",x"c1"),
  2947 => (x"02",x"9c",x"74",x"87"),
  2948 => (x"49",x"73",x"87",x"d8"),
  2949 => (x"99",x"c0",x"c0",x"c2"),
  2950 => (x"87",x"c3",x"c0",x"02"),
  2951 => (x"6d",x"2b",x"b7",x"d0"),
  2952 => (x"ff",x"ff",x"fd",x"48"),
  2953 => (x"c0",x"7d",x"70",x"98"),
  2954 => (x"d6",x"c4",x"87",x"f8"),
  2955 => (x"c0",x"02",x"bf",x"fc"),
  2956 => (x"48",x"73",x"87",x"f0"),
  2957 => (x"c8",x"28",x"b7",x"d0"),
  2958 => (x"98",x"70",x"58",x"a6"),
  2959 => (x"87",x"e2",x"c0",x"02"),
  2960 => (x"bf",x"c0",x"d7",x"c4"),
  2961 => (x"c0",x"e0",x"c0",x"49"),
  2962 => (x"ca",x"c0",x"02",x"99"),
  2963 => (x"c0",x"49",x"70",x"87"),
  2964 => (x"02",x"99",x"c0",x"e0"),
  2965 => (x"6d",x"87",x"cb",x"c0"),
  2966 => (x"c0",x"c0",x"c2",x"48"),
  2967 => (x"c4",x"7d",x"70",x"b0"),
  2968 => (x"49",x"73",x"4b",x"66"),
  2969 => (x"99",x"c0",x"c0",x"c8"),
  2970 => (x"87",x"c9",x"c2",x"02"),
  2971 => (x"bf",x"c0",x"d7",x"c4"),
  2972 => (x"9a",x"c0",x"cc",x"4a"),
  2973 => (x"87",x"cf",x"c0",x"02"),
  2974 => (x"02",x"8a",x"c0",x"c4"),
  2975 => (x"8a",x"87",x"d8",x"c0"),
  2976 => (x"87",x"fa",x"c0",x"02"),
  2977 => (x"73",x"87",x"df",x"c1"),
  2978 => (x"99",x"ff",x"c3",x"49"),
  2979 => (x"ef",x"c3",x"91",x"c2"),
  2980 => (x"4b",x"11",x"81",x"fc"),
  2981 => (x"73",x"87",x"de",x"c1"),
  2982 => (x"99",x"ff",x"c3",x"49"),
  2983 => (x"ef",x"c3",x"91",x"c2"),
  2984 => (x"81",x"c1",x"81",x"fc"),
  2985 => (x"9c",x"74",x"4b",x"11"),
  2986 => (x"87",x"c9",x"c0",x"02"),
  2987 => (x"48",x"a6",x"e0",x"c0"),
  2988 => (x"c0",x"c1",x"78",x"d2"),
  2989 => (x"48",x"a6",x"dc",x"87"),
  2990 => (x"c0",x"78",x"d2",x"c4"),
  2991 => (x"49",x"73",x"87",x"f7"),
  2992 => (x"c2",x"99",x"ff",x"c3"),
  2993 => (x"fc",x"ef",x"c3",x"91"),
  2994 => (x"11",x"81",x"c1",x"81"),
  2995 => (x"02",x"9c",x"74",x"4b"),
  2996 => (x"c0",x"87",x"ca",x"c0"),
  2997 => (x"c1",x"48",x"a6",x"e0"),
  2998 => (x"d8",x"c0",x"78",x"d9"),
  2999 => (x"48",x"a6",x"dc",x"87"),
  3000 => (x"c0",x"78",x"d9",x"c5"),
  3001 => (x"49",x"73",x"87",x"cf"),
  3002 => (x"c2",x"99",x"ff",x"c3"),
  3003 => (x"fc",x"ef",x"c3",x"91"),
  3004 => (x"11",x"81",x"c1",x"81"),
  3005 => (x"02",x"9c",x"74",x"4b"),
  3006 => (x"73",x"87",x"dc",x"c0"),
  3007 => (x"c7",x"b9",x"ff",x"49"),
  3008 => (x"71",x"99",x"c0",x"fc"),
  3009 => (x"c0",x"d7",x"c4",x"48"),
  3010 => (x"d7",x"c4",x"98",x"bf"),
  3011 => (x"ff",x"c3",x"58",x"c4"),
  3012 => (x"b3",x"c0",x"c4",x"9b"),
  3013 => (x"73",x"87",x"d4",x"c0"),
  3014 => (x"c0",x"fc",x"c7",x"49"),
  3015 => (x"c4",x"48",x"71",x"99"),
  3016 => (x"b0",x"bf",x"c0",x"d7"),
  3017 => (x"58",x"c4",x"d7",x"c4"),
  3018 => (x"dc",x"9b",x"ff",x"c3"),
  3019 => (x"ca",x"c0",x"02",x"66"),
  3020 => (x"d6",x"c4",x"1e",x"87"),
  3021 => (x"fb",x"f1",x"49",x"f4"),
  3022 => (x"73",x"86",x"c4",x"87"),
  3023 => (x"f4",x"d6",x"c4",x"1e"),
  3024 => (x"87",x"f0",x"f1",x"49"),
  3025 => (x"e0",x"c0",x"86",x"c4"),
  3026 => (x"ca",x"c0",x"02",x"66"),
  3027 => (x"d6",x"c4",x"1e",x"87"),
  3028 => (x"df",x"f1",x"49",x"f4"),
  3029 => (x"d4",x"86",x"c4",x"87"),
  3030 => (x"30",x"c1",x"48",x"66"),
  3031 => (x"6e",x"58",x"a6",x"d8"),
  3032 => (x"70",x"30",x"c1",x"48"),
  3033 => (x"48",x"66",x"d8",x"7e"),
  3034 => (x"a6",x"dc",x"80",x"c1"),
  3035 => (x"b7",x"e0",x"c0",x"58"),
  3036 => (x"f7",x"f8",x"04",x"a8"),
  3037 => (x"4c",x"66",x"d0",x"87"),
  3038 => (x"b7",x"c2",x"84",x"c1"),
  3039 => (x"e2",x"f7",x"04",x"ac"),
  3040 => (x"f8",x"d6",x"c4",x"87"),
  3041 => (x"78",x"66",x"c8",x"48"),
  3042 => (x"26",x"8e",x"dc",x"ff"),
  3043 => (x"26",x"4c",x"26",x"4d"),
  3044 => (x"00",x"4f",x"26",x"4b"),
  3045 => (x"00",x"00",x"00",x"00"),
  3046 => (x"72",x"4a",x"c0",x"1e"),
  3047 => (x"c4",x"91",x"c4",x"49"),
  3048 => (x"ff",x"81",x"c4",x"d7"),
  3049 => (x"c6",x"82",x"c1",x"79"),
  3050 => (x"ee",x"04",x"aa",x"b7"),
  3051 => (x"f8",x"d6",x"c4",x"87"),
  3052 => (x"40",x"40",x"c0",x"48"),
  3053 => (x"0e",x"4f",x"26",x"78"),
  3054 => (x"0e",x"5c",x"5b",x"5e"),
  3055 => (x"d4",x"ff",x"4a",x"71"),
  3056 => (x"4b",x"66",x"cc",x"4c"),
  3057 => (x"c8",x"48",x"d0",x"ff"),
  3058 => (x"7c",x"c2",x"78",x"c5"),
  3059 => (x"8b",x"c1",x"49",x"73"),
  3060 => (x"cd",x"02",x"99",x"71"),
  3061 => (x"12",x"7c",x"12",x"87"),
  3062 => (x"c1",x"49",x"73",x"7c"),
  3063 => (x"05",x"99",x"71",x"8b"),
  3064 => (x"d0",x"ff",x"87",x"f3"),
  3065 => (x"26",x"78",x"c4",x"48"),
  3066 => (x"26",x"4b",x"26",x"4c"),
  3067 => (x"4a",x"71",x"1e",x"4f"),
  3068 => (x"c8",x"48",x"d0",x"ff"),
  3069 => (x"d4",x"ff",x"78",x"c5"),
  3070 => (x"c8",x"78",x"c3",x"48"),
  3071 => (x"49",x"72",x"1e",x"c0"),
  3072 => (x"87",x"e3",x"c5",x"fd"),
  3073 => (x"c4",x"48",x"d0",x"ff"),
  3074 => (x"26",x"8e",x"fc",x"78"),
  3075 => (x"d0",x"ff",x"1e",x"4f"),
  3076 => (x"78",x"c5",x"c8",x"48"),
  3077 => (x"c6",x"48",x"d4",x"ff"),
  3078 => (x"ff",x"48",x"71",x"78"),
  3079 => (x"ff",x"78",x"08",x"d4"),
  3080 => (x"78",x"c4",x"48",x"d0"),
  3081 => (x"ff",x"1e",x"4f",x"26"),
  3082 => (x"c5",x"c8",x"48",x"d0"),
  3083 => (x"48",x"d4",x"ff",x"78"),
  3084 => (x"d0",x"ff",x"78",x"ca"),
  3085 => (x"26",x"78",x"c4",x"48"),
  3086 => (x"5b",x"5e",x"0e",x"4f"),
  3087 => (x"ff",x"0e",x"5d",x"5c"),
  3088 => (x"7e",x"71",x"86",x"d4"),
  3089 => (x"81",x"ca",x"49",x"6e"),
  3090 => (x"48",x"49",x"69",x"97"),
  3091 => (x"d4",x"28",x"b7",x"c5"),
  3092 => (x"49",x"6e",x"58",x"a6"),
  3093 => (x"69",x"97",x"81",x"c1"),
  3094 => (x"b7",x"c5",x"48",x"49"),
  3095 => (x"58",x"a6",x"d8",x"28"),
  3096 => (x"48",x"bf",x"97",x"6e"),
  3097 => (x"df",x"58",x"a6",x"dc"),
  3098 => (x"c0",x"c0",x"d0",x"99"),
  3099 => (x"c2",x"4a",x"6e",x"91"),
  3100 => (x"c0",x"48",x"12",x"82"),
  3101 => (x"70",x"58",x"a6",x"e0"),
  3102 => (x"92",x"c0",x"c4",x"4a"),
  3103 => (x"6e",x"49",x"a1",x"72"),
  3104 => (x"12",x"82",x"c3",x"4a"),
  3105 => (x"a6",x"e4",x"c0",x"48"),
  3106 => (x"c0",x"81",x"70",x"58"),
  3107 => (x"6e",x"59",x"a6",x"e8"),
  3108 => (x"c8",x"80",x"c4",x"48"),
  3109 => (x"66",x"c4",x"58",x"a6"),
  3110 => (x"9c",x"4c",x"bf",x"97"),
  3111 => (x"c4",x"87",x"c3",x"05"),
  3112 => (x"66",x"d0",x"4c",x"c0"),
  3113 => (x"a8",x"b7",x"c2",x"48"),
  3114 => (x"87",x"f1",x"cf",x"03"),
  3115 => (x"c1",x"49",x"66",x"d0"),
  3116 => (x"d4",x"c4",x"91",x"c8"),
  3117 => (x"80",x"71",x"48",x"e0"),
  3118 => (x"cc",x"58",x"a6",x"d0"),
  3119 => (x"80",x"c8",x"48",x"66"),
  3120 => (x"c8",x"58",x"a6",x"cc"),
  3121 => (x"cf",x"02",x"bf",x"66"),
  3122 => (x"c9",x"48",x"87",x"d3"),
  3123 => (x"a6",x"ec",x"c0",x"28"),
  3124 => (x"02",x"66",x"d8",x"58"),
  3125 => (x"4d",x"87",x"e3",x"c2"),
  3126 => (x"c3",x"02",x"8d",x"c3"),
  3127 => (x"8d",x"c1",x"87",x"c3"),
  3128 => (x"87",x"d6",x"c2",x"02"),
  3129 => (x"c4",x"02",x"8d",x"c4"),
  3130 => (x"8d",x"c2",x"87",x"cf"),
  3131 => (x"87",x"d6",x"c7",x"02"),
  3132 => (x"ca",x"02",x"8d",x"c8"),
  3133 => (x"02",x"8d",x"87",x"e5"),
  3134 => (x"cb",x"87",x"e6",x"cc"),
  3135 => (x"87",x"cf",x"02",x"8d"),
  3136 => (x"c3",x"02",x"8d",x"c3"),
  3137 => (x"8d",x"c2",x"87",x"f3"),
  3138 => (x"87",x"fa",x"c6",x"02"),
  3139 => (x"d4",x"87",x"fc",x"cd"),
  3140 => (x"d3",x"c1",x"05",x"66"),
  3141 => (x"d0",x"ff",x"c3",x"87"),
  3142 => (x"c8",x"4a",x"c0",x"4b"),
  3143 => (x"fe",x"fc",x"49",x"c0"),
  3144 => (x"e8",x"c0",x"87",x"f0"),
  3145 => (x"89",x"c1",x"49",x"66"),
  3146 => (x"2a",x"d8",x"4a",x"71"),
  3147 => (x"97",x"d4",x"ff",x"c3"),
  3148 => (x"d0",x"4a",x"71",x"5a"),
  3149 => (x"d5",x"ff",x"c3",x"2a"),
  3150 => (x"4a",x"71",x"5a",x"97"),
  3151 => (x"ff",x"c3",x"2a",x"c8"),
  3152 => (x"c3",x"5a",x"97",x"d6"),
  3153 => (x"59",x"97",x"d7",x"ff"),
  3154 => (x"c2",x"80",x"c3",x"48"),
  3155 => (x"f9",x"1e",x"c4",x"50"),
  3156 => (x"e2",x"f9",x"49",x"a0"),
  3157 => (x"c0",x"86",x"c4",x"87"),
  3158 => (x"87",x"f1",x"fa",x"49"),
  3159 => (x"49",x"e0",x"d3",x"c3"),
  3160 => (x"c0",x"81",x"66",x"d0"),
  3161 => (x"87",x"f8",x"cc",x"51"),
  3162 => (x"e0",x"fa",x"49",x"c2"),
  3163 => (x"e0",x"d3",x"c3",x"87"),
  3164 => (x"81",x"66",x"d0",x"49"),
  3165 => (x"cc",x"51",x"e5",x"c0"),
  3166 => (x"66",x"d4",x"87",x"e6"),
  3167 => (x"c3",x"87",x"d0",x"05"),
  3168 => (x"d0",x"49",x"e0",x"d3"),
  3169 => (x"51",x"c0",x"81",x"66"),
  3170 => (x"87",x"c1",x"fa",x"49"),
  3171 => (x"c3",x"87",x"d1",x"cc"),
  3172 => (x"d0",x"49",x"e0",x"d3"),
  3173 => (x"e5",x"c0",x"81",x"66"),
  3174 => (x"f9",x"49",x"c2",x"51"),
  3175 => (x"ff",x"cb",x"87",x"ef"),
  3176 => (x"02",x"66",x"d4",x"87"),
  3177 => (x"c3",x"87",x"ca",x"c0"),
  3178 => (x"d0",x"49",x"e0",x"d3"),
  3179 => (x"e5",x"c0",x"81",x"66"),
  3180 => (x"d0",x"ff",x"c3",x"51"),
  3181 => (x"c8",x"4a",x"c0",x"4b"),
  3182 => (x"fc",x"fc",x"49",x"c0"),
  3183 => (x"ff",x"c3",x"87",x"d4"),
  3184 => (x"50",x"cb",x"48",x"d7"),
  3185 => (x"48",x"e0",x"d3",x"c3"),
  3186 => (x"70",x"80",x"66",x"d0"),
  3187 => (x"bf",x"97",x"6e",x"7e"),
  3188 => (x"c0",x"02",x"99",x"49"),
  3189 => (x"ff",x"c3",x"87",x"cc"),
  3190 => (x"50",x"c5",x"48",x"d2"),
  3191 => (x"97",x"6e",x"80",x"c9"),
  3192 => (x"1e",x"c9",x"50",x"bf"),
  3193 => (x"49",x"d0",x"ff",x"c3"),
  3194 => (x"c4",x"87",x"cc",x"f7"),
  3195 => (x"f8",x"49",x"c0",x"86"),
  3196 => (x"48",x"6e",x"87",x"db"),
  3197 => (x"e7",x"ca",x"50",x"c0"),
  3198 => (x"05",x"66",x"d4",x"87"),
  3199 => (x"d8",x"87",x"f5",x"c2"),
  3200 => (x"e8",x"c0",x"48",x"66"),
  3201 => (x"c0",x"c1",x"05",x"a8"),
  3202 => (x"49",x"66",x"dc",x"87"),
  3203 => (x"c0",x"c0",x"c0",x"c1"),
  3204 => (x"e0",x"c0",x"91",x"c0"),
  3205 => (x"c0",x"d0",x"4a",x"66"),
  3206 => (x"a1",x"72",x"92",x"c0"),
  3207 => (x"97",x"66",x"c4",x"49"),
  3208 => (x"c0",x"c4",x"4a",x"bf"),
  3209 => (x"49",x"a1",x"72",x"92"),
  3210 => (x"82",x"c5",x"4a",x"6e"),
  3211 => (x"c0",x"4a",x"6a",x"97"),
  3212 => (x"72",x"48",x"a6",x"e4"),
  3213 => (x"49",x"6e",x"78",x"a1"),
  3214 => (x"69",x"97",x"81",x"c7"),
  3215 => (x"91",x"c0",x"c4",x"49"),
  3216 => (x"82",x"c8",x"4a",x"6e"),
  3217 => (x"a1",x"4a",x"6a",x"97"),
  3218 => (x"c0",x"49",x"74",x"4c"),
  3219 => (x"c0",x"81",x"66",x"e4"),
  3220 => (x"01",x"a9",x"66",x"e8"),
  3221 => (x"c0",x"87",x"cb",x"c1"),
  3222 => (x"c9",x"49",x"66",x"e4"),
  3223 => (x"d0",x"1e",x"71",x"31"),
  3224 => (x"e4",x"fd",x"49",x"66"),
  3225 => (x"86",x"c4",x"87",x"e5"),
  3226 => (x"8c",x"c1",x"49",x"74"),
  3227 => (x"c0",x"02",x"99",x"71"),
  3228 => (x"66",x"cc",x"87",x"df"),
  3229 => (x"75",x"1e",x"c0",x"4d"),
  3230 => (x"f4",x"de",x"fd",x"49"),
  3231 => (x"75",x"1e",x"c1",x"87"),
  3232 => (x"d1",x"dd",x"fd",x"49"),
  3233 => (x"74",x"86",x"c8",x"87"),
  3234 => (x"71",x"8c",x"c1",x"49"),
  3235 => (x"e4",x"ff",x"05",x"99"),
  3236 => (x"f5",x"49",x"c0",x"87"),
  3237 => (x"d3",x"c3",x"87",x"f7"),
  3238 => (x"66",x"d0",x"49",x"e0"),
  3239 => (x"c7",x"51",x"c0",x"81"),
  3240 => (x"49",x"c2",x"87",x"fe"),
  3241 => (x"c3",x"87",x"e6",x"f5"),
  3242 => (x"d0",x"49",x"e0",x"d3"),
  3243 => (x"e1",x"c0",x"81",x"66"),
  3244 => (x"87",x"ec",x"c7",x"51"),
  3245 => (x"d4",x"f5",x"49",x"c2"),
  3246 => (x"e0",x"d3",x"c3",x"87"),
  3247 => (x"81",x"66",x"d0",x"49"),
  3248 => (x"c7",x"51",x"e5",x"c0"),
  3249 => (x"66",x"d4",x"87",x"da"),
  3250 => (x"87",x"fd",x"c2",x"05"),
  3251 => (x"c0",x"48",x"66",x"d8"),
  3252 => (x"c1",x"05",x"a8",x"ea"),
  3253 => (x"66",x"dc",x"87",x"c0"),
  3254 => (x"c0",x"c0",x"c1",x"49"),
  3255 => (x"c0",x"91",x"c0",x"c0"),
  3256 => (x"d0",x"4a",x"66",x"e0"),
  3257 => (x"72",x"92",x"c0",x"c0"),
  3258 => (x"66",x"c4",x"49",x"a1"),
  3259 => (x"c4",x"4a",x"bf",x"97"),
  3260 => (x"a1",x"72",x"92",x"c0"),
  3261 => (x"c5",x"4a",x"6e",x"49"),
  3262 => (x"4a",x"6a",x"97",x"82"),
  3263 => (x"48",x"a6",x"e4",x"c0"),
  3264 => (x"6e",x"78",x"a1",x"72"),
  3265 => (x"97",x"81",x"c7",x"49"),
  3266 => (x"c0",x"c4",x"49",x"69"),
  3267 => (x"c8",x"4a",x"6e",x"91"),
  3268 => (x"4a",x"6a",x"97",x"82"),
  3269 => (x"49",x"74",x"4c",x"a1"),
  3270 => (x"81",x"66",x"e4",x"c0"),
  3271 => (x"a9",x"66",x"e8",x"c0"),
  3272 => (x"87",x"d3",x"c1",x"01"),
  3273 => (x"c0",x"02",x"9c",x"74"),
  3274 => (x"66",x"cc",x"87",x"fc"),
  3275 => (x"66",x"e4",x"c0",x"4d"),
  3276 => (x"71",x"31",x"c9",x"49"),
  3277 => (x"fd",x"49",x"75",x"1e"),
  3278 => (x"c3",x"87",x"d0",x"e1"),
  3279 => (x"f2",x"49",x"d0",x"ff"),
  3280 => (x"ff",x"c3",x"87",x"eb"),
  3281 => (x"49",x"75",x"1e",x"d0"),
  3282 => (x"87",x"f4",x"dc",x"fd"),
  3283 => (x"49",x"75",x"1e",x"c1"),
  3284 => (x"87",x"c2",x"da",x"fd"),
  3285 => (x"e4",x"c0",x"86",x"cc"),
  3286 => (x"80",x"c1",x"48",x"66"),
  3287 => (x"58",x"a6",x"e8",x"c0"),
  3288 => (x"ff",x"05",x"8c",x"c1"),
  3289 => (x"49",x"c0",x"87",x"c7"),
  3290 => (x"c3",x"87",x"e2",x"f2"),
  3291 => (x"d0",x"49",x"e0",x"d3"),
  3292 => (x"51",x"c0",x"81",x"66"),
  3293 => (x"c2",x"87",x"e9",x"c4"),
  3294 => (x"87",x"d1",x"f2",x"49"),
  3295 => (x"49",x"e0",x"d3",x"c3"),
  3296 => (x"c0",x"81",x"66",x"d0"),
  3297 => (x"d7",x"c4",x"51",x"e1"),
  3298 => (x"f1",x"49",x"c2",x"87"),
  3299 => (x"d3",x"c3",x"87",x"ff"),
  3300 => (x"66",x"d0",x"49",x"e0"),
  3301 => (x"51",x"e5",x"c0",x"81"),
  3302 => (x"c3",x"87",x"c5",x"c4"),
  3303 => (x"c0",x"4b",x"d0",x"ff"),
  3304 => (x"49",x"c0",x"c8",x"4a"),
  3305 => (x"87",x"ea",x"f4",x"fc"),
  3306 => (x"48",x"d2",x"ff",x"c3"),
  3307 => (x"49",x"74",x"50",x"c2"),
  3308 => (x"ff",x"c3",x"89",x"c5"),
  3309 => (x"c3",x"59",x"97",x"d8"),
  3310 => (x"c3",x"48",x"ec",x"d2"),
  3311 => (x"20",x"49",x"d8",x"ff"),
  3312 => (x"c3",x"41",x"20",x"41"),
  3313 => (x"c3",x"48",x"f8",x"d2"),
  3314 => (x"20",x"49",x"e0",x"ff"),
  3315 => (x"20",x"41",x"20",x"41"),
  3316 => (x"d0",x"41",x"20",x"41"),
  3317 => (x"f0",x"c0",x"49",x"66"),
  3318 => (x"f2",x"ff",x"c3",x"81"),
  3319 => (x"d3",x"c3",x"59",x"97"),
  3320 => (x"ff",x"c3",x"48",x"cc"),
  3321 => (x"41",x"20",x"49",x"f0"),
  3322 => (x"48",x"d4",x"d3",x"c3"),
  3323 => (x"49",x"f4",x"ff",x"c3"),
  3324 => (x"41",x"20",x"41",x"20"),
  3325 => (x"c0",x"02",x"66",x"d4"),
  3326 => (x"ff",x"c3",x"87",x"c7"),
  3327 => (x"ff",x"c1",x"48",x"d0"),
  3328 => (x"c1",x"49",x"74",x"50"),
  3329 => (x"c3",x"1e",x"71",x"29"),
  3330 => (x"ee",x"49",x"d0",x"ff"),
  3331 => (x"86",x"c4",x"87",x"e9"),
  3332 => (x"f8",x"ef",x"49",x"c0"),
  3333 => (x"e0",x"d3",x"c3",x"87"),
  3334 => (x"81",x"66",x"d0",x"49"),
  3335 => (x"ff",x"c1",x"51",x"c0"),
  3336 => (x"05",x"66",x"d4",x"87"),
  3337 => (x"c3",x"87",x"d2",x"c1"),
  3338 => (x"c0",x"4b",x"d0",x"ff"),
  3339 => (x"49",x"c0",x"c8",x"4a"),
  3340 => (x"87",x"de",x"f2",x"fc"),
  3341 => (x"48",x"d3",x"ff",x"c3"),
  3342 => (x"e8",x"c0",x"50",x"c8"),
  3343 => (x"29",x"d0",x"49",x"66"),
  3344 => (x"97",x"d9",x"ff",x"c3"),
  3345 => (x"66",x"e8",x"c0",x"59"),
  3346 => (x"c3",x"29",x"c8",x"49"),
  3347 => (x"59",x"97",x"da",x"ff"),
  3348 => (x"c0",x"80",x"c1",x"48"),
  3349 => (x"c2",x"50",x"66",x"e8"),
  3350 => (x"49",x"74",x"50",x"80"),
  3351 => (x"1e",x"71",x"29",x"c1"),
  3352 => (x"ed",x"49",x"a0",x"f5"),
  3353 => (x"86",x"c4",x"87",x"d1"),
  3354 => (x"e0",x"ee",x"49",x"c0"),
  3355 => (x"e0",x"d3",x"c3",x"87"),
  3356 => (x"81",x"66",x"d0",x"49"),
  3357 => (x"e7",x"c0",x"51",x"c0"),
  3358 => (x"e0",x"d3",x"c3",x"87"),
  3359 => (x"81",x"66",x"d0",x"49"),
  3360 => (x"c2",x"51",x"e5",x"c0"),
  3361 => (x"87",x"c5",x"ee",x"49"),
  3362 => (x"c3",x"87",x"d5",x"c0"),
  3363 => (x"d0",x"49",x"e0",x"d3"),
  3364 => (x"e0",x"c0",x"81",x"66"),
  3365 => (x"ed",x"49",x"c2",x"51"),
  3366 => (x"c3",x"c0",x"87",x"f3"),
  3367 => (x"87",x"c6",x"ee",x"87"),
  3368 => (x"26",x"8e",x"d4",x"ff"),
  3369 => (x"26",x"4c",x"26",x"4d"),
  3370 => (x"00",x"4f",x"26",x"4b"),
  3371 => (x"34",x"36",x"43",x"54"),
  3372 => (x"20",x"20",x"20",x"20"),
  3373 => (x"00",x"00",x"00",x"00"),
  3374 => (x"69",x"4d",x"65",x"44"),
  3375 => (x"66",x"69",x"54",x"53"),
  3376 => (x"44",x"48",x"20",x"79"),
  3377 => (x"20",x"30",x"20",x"44"),
  3378 => (x"00",x"00",x"00",x"00"),
  3379 => (x"20",x"32",x"33",x"38"),
  3380 => (x"00",x"00",x"00",x"00"),
  3381 => (x"32",x"31",x"30",x"32"),
  3382 => (x"39",x"32",x"39",x"30"),
  3383 => (x"00",x"00",x"00",x"09"),
  3384 => (x"73",x"1e",x"00",x"00"),
  3385 => (x"ff",x"86",x"e0",x"1e"),
  3386 => (x"c5",x"c8",x"48",x"d0"),
  3387 => (x"48",x"d4",x"ff",x"78"),
  3388 => (x"1e",x"d0",x"78",x"c5"),
  3389 => (x"49",x"4b",x"a6",x"c4"),
  3390 => (x"87",x"eb",x"f1",x"fc"),
  3391 => (x"d0",x"ff",x"86",x"c4"),
  3392 => (x"ca",x"78",x"c4",x"48"),
  3393 => (x"c1",x"49",x"66",x"97"),
  3394 => (x"87",x"c5",x"02",x"99"),
  3395 => (x"e8",x"ec",x"49",x"73"),
  3396 => (x"26",x"8e",x"e0",x"87"),
  3397 => (x"1e",x"4f",x"26",x"4b"),
  3398 => (x"c4",x"4a",x"d4",x"ff"),
  3399 => (x"c4",x"48",x"f8",x"d7"),
  3400 => (x"78",x"bf",x"e4",x"d1"),
  3401 => (x"ff",x"7a",x"ff",x"c3"),
  3402 => (x"78",x"c5",x"48",x"d0"),
  3403 => (x"d1",x"c4",x"7a",x"c4"),
  3404 => (x"48",x"49",x"bf",x"e4"),
  3405 => (x"7a",x"70",x"28",x"d8"),
  3406 => (x"28",x"d0",x"48",x"71"),
  3407 => (x"48",x"71",x"7a",x"70"),
  3408 => (x"7a",x"70",x"28",x"c8"),
  3409 => (x"bf",x"e4",x"d1",x"c4"),
  3410 => (x"48",x"d0",x"ff",x"7a"),
  3411 => (x"4f",x"26",x"78",x"c4"),
  3412 => (x"c4",x"4a",x"c0",x"1e"),
  3413 => (x"02",x"bf",x"ec",x"d8"),
  3414 => (x"c4",x"49",x"87",x"ca"),
  3415 => (x"c1",x"48",x"ec",x"d8"),
  3416 => (x"4a",x"11",x"78",x"a1"),
  3417 => (x"c6",x"05",x"9a",x"72"),
  3418 => (x"ec",x"d8",x"c4",x"87"),
  3419 => (x"72",x"78",x"c0",x"48"),
  3420 => (x"1e",x"4f",x"26",x"48"),
  3421 => (x"48",x"ec",x"d8",x"c4"),
  3422 => (x"bf",x"c8",x"f4",x"c3"),
  3423 => (x"0e",x"4f",x"26",x"78"),
  3424 => (x"0e",x"5c",x"5b",x"5e"),
  3425 => (x"d0",x"ff",x"4a",x"71"),
  3426 => (x"4b",x"d4",x"ff",x"4c"),
  3427 => (x"d5",x"c1",x"7c",x"c5"),
  3428 => (x"7b",x"66",x"cc",x"7b"),
  3429 => (x"7c",x"c5",x"7c",x"c4"),
  3430 => (x"c1",x"7b",x"d3",x"c1"),
  3431 => (x"c8",x"7c",x"c4",x"7b"),
  3432 => (x"d4",x"c1",x"7c",x"c5"),
  3433 => (x"b7",x"49",x"c0",x"7b"),
  3434 => (x"87",x"ca",x"06",x"aa"),
  3435 => (x"81",x"c1",x"7b",x"c0"),
  3436 => (x"04",x"a9",x"b7",x"72"),
  3437 => (x"7c",x"c4",x"87",x"f6"),
  3438 => (x"d3",x"c1",x"7c",x"c5"),
  3439 => (x"c4",x"7b",x"c0",x"7b"),
  3440 => (x"26",x"4c",x"26",x"7c"),
  3441 => (x"1e",x"4f",x"26",x"4b"),
  3442 => (x"4b",x"71",x"1e",x"73"),
  3443 => (x"97",x"e0",x"f3",x"c1"),
  3444 => (x"b7",x"c2",x"49",x"bf"),
  3445 => (x"f3",x"c0",x"03",x"a9"),
  3446 => (x"c4",x"1e",x"73",x"87"),
  3447 => (x"fd",x"49",x"cc",x"cc"),
  3448 => (x"c4",x"87",x"d0",x"cb"),
  3449 => (x"02",x"98",x"70",x"86"),
  3450 => (x"c4",x"87",x"e1",x"c0"),
  3451 => (x"4a",x"bf",x"d4",x"cc"),
  3452 => (x"c0",x"c3",x"2a",x"ca"),
  3453 => (x"87",x"ce",x"02",x"8a"),
  3454 => (x"05",x"8a",x"c0",x"c1"),
  3455 => (x"f3",x"c1",x"87",x"ce"),
  3456 => (x"50",x"c0",x"48",x"e0"),
  3457 => (x"f3",x"c1",x"87",x"c6"),
  3458 => (x"50",x"c1",x"48",x"e0"),
  3459 => (x"4f",x"26",x"4b",x"26"),
  3460 => (x"71",x"1e",x"73",x"1e"),
  3461 => (x"c6",x"02",x"9a",x"4a"),
  3462 => (x"c4",x"dd",x"c3",x"87"),
  3463 => (x"c3",x"78",x"c0",x"48"),
  3464 => (x"49",x"bf",x"c0",x"dd"),
  3465 => (x"87",x"c0",x"ce",x"ff"),
  3466 => (x"c4",x"02",x"98",x"70"),
  3467 => (x"49",x"d4",x"87",x"cd"),
  3468 => (x"87",x"e8",x"cd",x"ff"),
  3469 => (x"58",x"c4",x"dd",x"c3"),
  3470 => (x"bf",x"c4",x"dd",x"c3"),
  3471 => (x"87",x"fb",x"c0",x"05"),
  3472 => (x"49",x"d0",x"d1",x"c4"),
  3473 => (x"87",x"ce",x"df",x"fe"),
  3474 => (x"04",x"a8",x"b7",x"c0"),
  3475 => (x"d1",x"c4",x"87",x"ce"),
  3476 => (x"df",x"fe",x"49",x"d0"),
  3477 => (x"b7",x"c0",x"87",x"c0"),
  3478 => (x"87",x"f2",x"03",x"a8"),
  3479 => (x"bf",x"c4",x"dd",x"c3"),
  3480 => (x"c4",x"dd",x"c3",x"49"),
  3481 => (x"78",x"a1",x"c1",x"48"),
  3482 => (x"81",x"cc",x"f4",x"c3"),
  3483 => (x"dd",x"c3",x"48",x"11"),
  3484 => (x"dd",x"c3",x"58",x"cc"),
  3485 => (x"78",x"c0",x"48",x"cc"),
  3486 => (x"c3",x"87",x"c0",x"c3"),
  3487 => (x"02",x"bf",x"cc",x"dd"),
  3488 => (x"c4",x"87",x"f5",x"c1"),
  3489 => (x"fe",x"49",x"d0",x"d1"),
  3490 => (x"c0",x"87",x"cb",x"de"),
  3491 => (x"cd",x"04",x"a8",x"b7"),
  3492 => (x"cc",x"dd",x"c3",x"87"),
  3493 => (x"88",x"c1",x"48",x"bf"),
  3494 => (x"58",x"d0",x"dd",x"c3"),
  3495 => (x"d6",x"c4",x"87",x"dd"),
  3496 => (x"ff",x"49",x"bf",x"f0"),
  3497 => (x"70",x"87",x"c1",x"cc"),
  3498 => (x"ce",x"c0",x"02",x"98"),
  3499 => (x"d0",x"d1",x"c4",x"87"),
  3500 => (x"d6",x"db",x"fe",x"49"),
  3501 => (x"c4",x"dd",x"c3",x"87"),
  3502 => (x"c3",x"78",x"c0",x"48"),
  3503 => (x"05",x"bf",x"c8",x"dd"),
  3504 => (x"c3",x"87",x"f8",x"c1"),
  3505 => (x"05",x"bf",x"cc",x"dd"),
  3506 => (x"c3",x"87",x"f0",x"c1"),
  3507 => (x"49",x"bf",x"c4",x"dd"),
  3508 => (x"48",x"c4",x"dd",x"c3"),
  3509 => (x"c3",x"78",x"a1",x"c1"),
  3510 => (x"11",x"81",x"cc",x"f4"),
  3511 => (x"c0",x"c2",x"49",x"4b"),
  3512 => (x"cc",x"c0",x"02",x"99"),
  3513 => (x"c1",x"48",x"73",x"87"),
  3514 => (x"dd",x"c3",x"98",x"ff"),
  3515 => (x"ca",x"c1",x"58",x"d0"),
  3516 => (x"cc",x"dd",x"c3",x"87"),
  3517 => (x"87",x"c3",x"c1",x"5b"),
  3518 => (x"bf",x"c8",x"dd",x"c3"),
  3519 => (x"87",x"fb",x"c0",x"02"),
  3520 => (x"bf",x"c4",x"dd",x"c3"),
  3521 => (x"c4",x"dd",x"c3",x"49"),
  3522 => (x"78",x"a1",x"c1",x"48"),
  3523 => (x"81",x"cc",x"f4",x"c3"),
  3524 => (x"1e",x"49",x"69",x"97"),
  3525 => (x"49",x"d0",x"d1",x"c4"),
  3526 => (x"87",x"c6",x"da",x"fe"),
  3527 => (x"dd",x"c3",x"86",x"c4"),
  3528 => (x"c1",x"48",x"bf",x"c8"),
  3529 => (x"cc",x"dd",x"c3",x"88"),
  3530 => (x"cc",x"dd",x"c3",x"58"),
  3531 => (x"c0",x"78",x"c1",x"48"),
  3532 => (x"ff",x"49",x"ec",x"f6"),
  3533 => (x"c4",x"87",x"e5",x"c9"),
  3534 => (x"26",x"58",x"f4",x"d6"),
  3535 => (x"00",x"4f",x"26",x"4b"),
  3536 => (x"00",x"00",x"00",x"00"),
  3537 => (x"00",x"00",x"00",x"00"),
  3538 => (x"00",x"00",x"00",x"00"),
  3539 => (x"00",x"00",x"00",x"00"),
  3540 => (x"71",x"1e",x"73",x"1e"),
  3541 => (x"fb",x"fd",x"49",x"4b"),
  3542 => (x"d1",x"c4",x"87",x"f0"),
  3543 => (x"02",x"bf",x"97",x"f8"),
  3544 => (x"1e",x"c3",x"87",x"cb"),
  3545 => (x"49",x"c0",x"c0",x"c4"),
  3546 => (x"c4",x"87",x"d4",x"f8"),
  3547 => (x"fd",x"49",x"73",x"86"),
  3548 => (x"26",x"87",x"d7",x"fb"),
  3549 => (x"1e",x"4f",x"26",x"4b"),
  3550 => (x"da",x"f6",x"1e",x"73"),
  3551 => (x"49",x"f4",x"c7",x"87"),
  3552 => (x"87",x"d8",x"c8",x"ff"),
  3553 => (x"ff",x"49",x"4b",x"70"),
  3554 => (x"70",x"87",x"dd",x"c8"),
  3555 => (x"87",x"cb",x"05",x"98"),
  3556 => (x"c8",x"ff",x"49",x"73"),
  3557 => (x"98",x"70",x"87",x"d2"),
  3558 => (x"26",x"87",x"f5",x"02"),
  3559 => (x"0e",x"4f",x"26",x"4b"),
  3560 => (x"5d",x"5c",x"5b",x"5e"),
  3561 => (x"71",x"86",x"f8",x"0e"),
  3562 => (x"fd",x"4d",x"c0",x"4b"),
  3563 => (x"70",x"87",x"ee",x"d4"),
  3564 => (x"02",x"9b",x"73",x"4c"),
  3565 => (x"c1",x"87",x"c2",x"c5"),
  3566 => (x"c1",x"48",x"e0",x"f3"),
  3567 => (x"c4",x"1e",x"73",x"50"),
  3568 => (x"fd",x"49",x"cc",x"cc"),
  3569 => (x"c4",x"87",x"ec",x"c3"),
  3570 => (x"02",x"98",x"70",x"86"),
  3571 => (x"c4",x"87",x"ff",x"c3"),
  3572 => (x"48",x"bf",x"e4",x"d1"),
  3573 => (x"d1",x"c4",x"b0",x"c1"),
  3574 => (x"fa",x"f4",x"58",x"e8"),
  3575 => (x"d0",x"ff",x"c3",x"87"),
  3576 => (x"cc",x"cc",x"c4",x"1e"),
  3577 => (x"c8",x"c9",x"fd",x"49"),
  3578 => (x"c3",x"86",x"c4",x"87"),
  3579 => (x"7e",x"bf",x"dc",x"ff"),
  3580 => (x"c3",x"48",x"a6",x"c4"),
  3581 => (x"78",x"bf",x"e0",x"ff"),
  3582 => (x"97",x"d0",x"ff",x"c3"),
  3583 => (x"a9",x"c1",x"49",x"bf"),
  3584 => (x"87",x"ca",x"c3",x"05"),
  3585 => (x"bf",x"d4",x"ff",x"c3"),
  3586 => (x"71",x"b1",x"c1",x"49"),
  3587 => (x"ff",x"cf",x"ff",x"48"),
  3588 => (x"e8",x"d1",x"c4",x"98"),
  3589 => (x"d1",x"ff",x"c3",x"58"),
  3590 => (x"c2",x"48",x"bf",x"97"),
  3591 => (x"c3",x"58",x"d0",x"e6"),
  3592 => (x"49",x"bf",x"d8",x"ff"),
  3593 => (x"87",x"f2",x"dd",x"fd"),
  3594 => (x"c0",x"02",x"98",x"70"),
  3595 => (x"ff",x"c3",x"87",x"e2"),
  3596 => (x"cc",x"c4",x"1e",x"d0"),
  3597 => (x"c7",x"fd",x"49",x"cc"),
  3598 => (x"ff",x"c3",x"87",x"f7"),
  3599 => (x"fd",x"49",x"bf",x"d8"),
  3600 => (x"c0",x"87",x"fb",x"d0"),
  3601 => (x"e4",x"ff",x"c3",x"1e"),
  3602 => (x"87",x"cc",x"c4",x"49"),
  3603 => (x"4d",x"70",x"86",x"c8"),
  3604 => (x"d0",x"fd",x"49",x"74"),
  3605 => (x"1e",x"73",x"87",x"e8"),
  3606 => (x"49",x"cc",x"cc",x"c4"),
  3607 => (x"87",x"d3",x"c1",x"fd"),
  3608 => (x"49",x"6e",x"86",x"c4"),
  3609 => (x"87",x"f2",x"dc",x"fd"),
  3610 => (x"c0",x"02",x"98",x"70"),
  3611 => (x"ff",x"c3",x"87",x"e1"),
  3612 => (x"cc",x"c4",x"1e",x"d0"),
  3613 => (x"c6",x"fd",x"49",x"cc"),
  3614 => (x"ff",x"c3",x"87",x"f7"),
  3615 => (x"fd",x"49",x"bf",x"dc"),
  3616 => (x"c0",x"87",x"fb",x"cf"),
  3617 => (x"ff",x"c3",x"1e",x"f2"),
  3618 => (x"cb",x"c3",x"49",x"f0"),
  3619 => (x"74",x"86",x"c8",x"87"),
  3620 => (x"e9",x"cf",x"fd",x"49"),
  3621 => (x"c4",x"1e",x"73",x"87"),
  3622 => (x"fd",x"49",x"cc",x"cc"),
  3623 => (x"c4",x"87",x"d4",x"c0"),
  3624 => (x"fd",x"49",x"66",x"86"),
  3625 => (x"70",x"87",x"f3",x"db"),
  3626 => (x"e1",x"c0",x"02",x"98"),
  3627 => (x"d0",x"ff",x"c3",x"87"),
  3628 => (x"cc",x"cc",x"c4",x"1e"),
  3629 => (x"f8",x"c5",x"fd",x"49"),
  3630 => (x"e0",x"ff",x"c3",x"87"),
  3631 => (x"ce",x"fd",x"49",x"bf"),
  3632 => (x"f3",x"c0",x"87",x"fc"),
  3633 => (x"fc",x"ff",x"c3",x"1e"),
  3634 => (x"87",x"cc",x"c2",x"49"),
  3635 => (x"1e",x"c2",x"86",x"c8"),
  3636 => (x"49",x"c0",x"c0",x"c4"),
  3637 => (x"c3",x"87",x"e8",x"f2"),
  3638 => (x"c0",x"c0",x"c4",x"1e"),
  3639 => (x"87",x"df",x"f2",x"49"),
  3640 => (x"d1",x"c4",x"86",x"c8"),
  3641 => (x"fe",x"48",x"bf",x"e4"),
  3642 => (x"e8",x"d1",x"c4",x"98"),
  3643 => (x"87",x"e7",x"f0",x"58"),
  3644 => (x"bf",x"cc",x"e6",x"c2"),
  3645 => (x"d2",x"f5",x"fe",x"49"),
  3646 => (x"f8",x"48",x"75",x"87"),
  3647 => (x"26",x"4d",x"26",x"8e"),
  3648 => (x"26",x"4b",x"26",x"4c"),
  3649 => (x"1e",x"73",x"1e",x"4f"),
  3650 => (x"49",x"ca",x"4b",x"71"),
  3651 => (x"87",x"fe",x"dc",x"fc"),
  3652 => (x"cc",x"c4",x"1e",x"73"),
  3653 => (x"fe",x"fc",x"49",x"cc"),
  3654 => (x"86",x"c4",x"87",x"d9"),
  3655 => (x"c0",x"02",x"98",x"70"),
  3656 => (x"d7",x"c4",x"87",x"f0"),
  3657 => (x"50",x"c1",x"48",x"f4"),
  3658 => (x"bf",x"cc",x"e6",x"c2"),
  3659 => (x"c4",x"80",x"c2",x"50"),
  3660 => (x"78",x"bf",x"e4",x"d1"),
  3661 => (x"50",x"c0",x"80",x"db"),
  3662 => (x"50",x"c0",x"80",x"cb"),
  3663 => (x"50",x"c0",x"80",x"cb"),
  3664 => (x"1e",x"a0",x"c8",x"ff"),
  3665 => (x"49",x"cc",x"cc",x"c4"),
  3666 => (x"87",x"f4",x"c4",x"fd"),
  3667 => (x"48",x"c1",x"86",x"c4"),
  3668 => (x"48",x"c0",x"87",x"c2"),
  3669 => (x"4f",x"26",x"4b",x"26"),
  3670 => (x"5c",x"5b",x"5e",x"0e"),
  3671 => (x"86",x"f4",x"0e",x"5d"),
  3672 => (x"7e",x"c0",x"4d",x"71"),
  3673 => (x"c0",x"48",x"66",x"dc"),
  3674 => (x"a6",x"cc",x"88",x"f0"),
  3675 => (x"02",x"66",x"dc",x"58"),
  3676 => (x"70",x"87",x"e6",x"c0"),
  3677 => (x"f3",x"c1",x"02",x"98"),
  3678 => (x"8c",x"c1",x"4c",x"87"),
  3679 => (x"87",x"ec",x"c1",x"02"),
  3680 => (x"d1",x"c2",x"02",x"8c"),
  3681 => (x"c2",x"02",x"8c",x"87"),
  3682 => (x"8c",x"d0",x"87",x"cc"),
  3683 => (x"87",x"e7",x"c4",x"02"),
  3684 => (x"c4",x"02",x"8c",x"c1"),
  3685 => (x"ef",x"c4",x"87",x"eb"),
  3686 => (x"02",x"9d",x"75",x"87"),
  3687 => (x"97",x"87",x"e9",x"c4"),
  3688 => (x"e3",x"c4",x"02",x"6d"),
  3689 => (x"c4",x"1e",x"c2",x"87"),
  3690 => (x"ef",x"49",x"c0",x"c0"),
  3691 => (x"86",x"c4",x"87",x"d1"),
  3692 => (x"4b",x"c8",x"d8",x"c4"),
  3693 => (x"49",x"cb",x"4a",x"75"),
  3694 => (x"87",x"c6",x"dc",x"fc"),
  3695 => (x"48",x"d3",x"d8",x"c4"),
  3696 => (x"cc",x"fd",x"50",x"c0"),
  3697 => (x"d8",x"c4",x"87",x"d7"),
  3698 => (x"d1",x"c4",x"58",x"c0"),
  3699 => (x"c1",x"48",x"bf",x"e4"),
  3700 => (x"e8",x"d1",x"c4",x"b0"),
  3701 => (x"87",x"ff",x"ec",x"58"),
  3702 => (x"49",x"c8",x"d8",x"c4"),
  3703 => (x"c4",x"87",x"e8",x"ef"),
  3704 => (x"fd",x"49",x"c8",x"d8"),
  3705 => (x"c1",x"87",x"de",x"e0"),
  3706 => (x"87",x"dc",x"c3",x"7e"),
  3707 => (x"c0",x"1e",x"66",x"c8"),
  3708 => (x"d7",x"c4",x"ff",x"49"),
  3709 => (x"49",x"66",x"cc",x"87"),
  3710 => (x"cc",x"87",x"fc",x"f5"),
  3711 => (x"49",x"75",x"1e",x"66"),
  3712 => (x"87",x"c8",x"c4",x"ff"),
  3713 => (x"49",x"66",x"86",x"c8"),
  3714 => (x"c4",x"91",x"c8",x"c1"),
  3715 => (x"c8",x"81",x"d0",x"d2"),
  3716 => (x"c2",x"7e",x"69",x"81"),
  3717 => (x"66",x"c8",x"87",x"f2"),
  3718 => (x"91",x"c8",x"c1",x"49"),
  3719 => (x"48",x"d0",x"d2",x"c4"),
  3720 => (x"7e",x"70",x"80",x"71"),
  3721 => (x"a6",x"80",x"c8",x"48"),
  3722 => (x"48",x"66",x"c4",x"58"),
  3723 => (x"9d",x"75",x"78",x"c0"),
  3724 => (x"87",x"e6",x"c0",x"02"),
  3725 => (x"cc",x"4c",x"66",x"c8"),
  3726 => (x"fc",x"d7",x"c4",x"94"),
  3727 => (x"75",x"4b",x"74",x"84"),
  3728 => (x"fc",x"49",x"cb",x"4a"),
  3729 => (x"cb",x"87",x"fb",x"d9"),
  3730 => (x"51",x"c0",x"49",x"a4"),
  3731 => (x"66",x"c4",x"1e",x"74"),
  3732 => (x"de",x"f9",x"fc",x"49"),
  3733 => (x"c0",x"86",x"c4",x"87"),
  3734 => (x"66",x"c8",x"87",x"cb"),
  3735 => (x"c4",x"91",x"cc",x"49"),
  3736 => (x"c0",x"81",x"fc",x"d7"),
  3737 => (x"f4",x"c9",x"fd",x"51"),
  3738 => (x"c8",x"4a",x"70",x"87"),
  3739 => (x"91",x"c4",x"49",x"66"),
  3740 => (x"81",x"f8",x"d7",x"c4"),
  3741 => (x"66",x"c4",x"79",x"72"),
  3742 => (x"da",x"c0",x"02",x"bf"),
  3743 => (x"49",x"66",x"c8",x"87"),
  3744 => (x"c0",x"d0",x"89",x"c2"),
  3745 => (x"70",x"30",x"71",x"48"),
  3746 => (x"e4",x"d1",x"c4",x"49"),
  3747 => (x"b0",x"71",x"48",x"bf"),
  3748 => (x"58",x"e8",x"d1",x"c4"),
  3749 => (x"c8",x"87",x"d9",x"c0"),
  3750 => (x"89",x"c2",x"49",x"66"),
  3751 => (x"71",x"48",x"c0",x"d0"),
  3752 => (x"ff",x"49",x"70",x"30"),
  3753 => (x"e4",x"d1",x"c4",x"b9"),
  3754 => (x"98",x"71",x"48",x"bf"),
  3755 => (x"58",x"e8",x"d1",x"c4"),
  3756 => (x"7e",x"bf",x"66",x"c4"),
  3757 => (x"75",x"87",x"d1",x"c0"),
  3758 => (x"87",x"e3",x"f3",x"49"),
  3759 => (x"c7",x"c0",x"7e",x"70"),
  3760 => (x"f8",x"49",x"75",x"87"),
  3761 => (x"7e",x"70",x"87",x"ff"),
  3762 => (x"bf",x"e4",x"d1",x"c4"),
  3763 => (x"c4",x"98",x"fe",x"48"),
  3764 => (x"e9",x"58",x"e8",x"d1"),
  3765 => (x"48",x"6e",x"87",x"c1"),
  3766 => (x"4d",x"26",x"8e",x"f4"),
  3767 => (x"4b",x"26",x"4c",x"26"),
  3768 => (x"73",x"1e",x"4f",x"26"),
  3769 => (x"e4",x"d1",x"c4",x"1e"),
  3770 => (x"c1",x"78",x"c1",x"48"),
  3771 => (x"c1",x"48",x"e0",x"f3"),
  3772 => (x"c4",x"c8",x"c1",x"50"),
  3773 => (x"e8",x"50",x"c0",x"48"),
  3774 => (x"1e",x"c3",x"87",x"dd"),
  3775 => (x"49",x"c0",x"c0",x"c4"),
  3776 => (x"c2",x"87",x"fc",x"e9"),
  3777 => (x"c0",x"c0",x"c4",x"1e"),
  3778 => (x"87",x"f3",x"e9",x"49"),
  3779 => (x"f4",x"c3",x"86",x"c8"),
  3780 => (x"f2",x"49",x"bf",x"e0"),
  3781 => (x"98",x"70",x"87",x"c9"),
  3782 => (x"87",x"ef",x"c1",x"05"),
  3783 => (x"c3",x"87",x"f8",x"e7"),
  3784 => (x"49",x"bf",x"dc",x"f4"),
  3785 => (x"c3",x"87",x"e0",x"ea"),
  3786 => (x"49",x"bf",x"dc",x"f4"),
  3787 => (x"87",x"d5",x"db",x"fd"),
  3788 => (x"bf",x"e4",x"d1",x"c4"),
  3789 => (x"c4",x"98",x"fe",x"48"),
  3790 => (x"e7",x"58",x"e8",x"d1"),
  3791 => (x"d0",x"c6",x"87",x"d9"),
  3792 => (x"d7",x"f9",x"fe",x"49"),
  3793 => (x"49",x"4b",x"70",x"87"),
  3794 => (x"87",x"dc",x"f9",x"fe"),
  3795 => (x"cc",x"05",x"98",x"70"),
  3796 => (x"fe",x"49",x"73",x"87"),
  3797 => (x"70",x"87",x"d1",x"f9"),
  3798 => (x"f4",x"ff",x"02",x"98"),
  3799 => (x"e4",x"d1",x"c4",x"87"),
  3800 => (x"b0",x"c1",x"48",x"bf"),
  3801 => (x"58",x"e8",x"d1",x"c4"),
  3802 => (x"c1",x"87",x"ec",x"e6"),
  3803 => (x"f8",x"fe",x"49",x"e4"),
  3804 => (x"4b",x"70",x"87",x"ea"),
  3805 => (x"ef",x"f8",x"fe",x"49"),
  3806 => (x"05",x"98",x"70",x"87"),
  3807 => (x"73",x"87",x"cc",x"c0"),
  3808 => (x"e3",x"f8",x"fe",x"49"),
  3809 => (x"02",x"98",x"70",x"87"),
  3810 => (x"c4",x"87",x"f4",x"ff"),
  3811 => (x"48",x"bf",x"e4",x"d1"),
  3812 => (x"d1",x"c4",x"98",x"fe"),
  3813 => (x"fe",x"e5",x"58",x"e8"),
  3814 => (x"fb",x"cf",x"ff",x"87"),
  3815 => (x"da",x"c7",x"fe",x"87"),
  3816 => (x"e9",x"49",x"c1",x"87"),
  3817 => (x"48",x"c0",x"87",x"ea"),
  3818 => (x"4f",x"26",x"4b",x"26"),
  3819 => (x"71",x"1e",x"73",x"1e"),
  3820 => (x"cf",x"c4",x"ff",x"4b"),
  3821 => (x"fe",x"49",x"73",x"87"),
  3822 => (x"26",x"87",x"d0",x"cf"),
  3823 => (x"0e",x"4f",x"26",x"4b"),
  3824 => (x"0e",x"5c",x"5b",x"5e"),
  3825 => (x"ff",x"c1",x"86",x"fc"),
  3826 => (x"4b",x"6e",x"4c",x"ff"),
  3827 => (x"ff",x"e8",x"49",x"c0"),
  3828 => (x"de",x"ed",x"fe",x"87"),
  3829 => (x"dc",x"f9",x"fe",x"87"),
  3830 => (x"87",x"c6",x"e4",x"87"),
  3831 => (x"99",x"74",x"49",x"73"),
  3832 => (x"99",x"71",x"83",x"c1"),
  3833 => (x"fd",x"87",x"e5",x"05"),
  3834 => (x"70",x"87",x"f9",x"ff"),
  3835 => (x"ee",x"d4",x"fe",x"49"),
  3836 => (x"87",x"d8",x"ff",x"87"),
  3837 => (x"4c",x"26",x"8e",x"fc"),
  3838 => (x"4f",x"26",x"4b",x"26"),
  3839 => (x"f5",x"f2",x"eb",x"f4"),
  3840 => (x"0c",x"04",x"06",x"05"),
  3841 => (x"0a",x"83",x"0b",x"03"),
  3842 => (x"00",x"00",x"00",x"66"),
  3843 => (x"00",x"da",x"00",x"5a"),
  3844 => (x"08",x"94",x"80",x"00"),
  3845 => (x"00",x"78",x"80",x"05"),
  3846 => (x"00",x"01",x"80",x"02"),
  3847 => (x"00",x"09",x"80",x"03"),
  3848 => (x"00",x"00",x"80",x"04"),
  3849 => (x"08",x"91",x"80",x"01"),
  3850 => (x"00",x"00",x"00",x"26"),
  3851 => (x"00",x"00",x"00",x"1d"),
  3852 => (x"00",x"00",x"00",x"1c"),
  3853 => (x"00",x"00",x"00",x"25"),
  3854 => (x"00",x"00",x"00",x"1a"),
  3855 => (x"00",x"00",x"00",x"1b"),
  3856 => (x"00",x"00",x"00",x"24"),
  3857 => (x"00",x"00",x"01",x"12"),
  3858 => (x"00",x"00",x"00",x"2e"),
  3859 => (x"00",x"00",x"00",x"2d"),
  3860 => (x"00",x"00",x"00",x"23"),
  3861 => (x"00",x"00",x"00",x"36"),
  3862 => (x"00",x"00",x"00",x"21"),
  3863 => (x"00",x"00",x"00",x"2b"),
  3864 => (x"00",x"00",x"00",x"2c"),
  3865 => (x"00",x"00",x"00",x"22"),
  3866 => (x"00",x"6c",x"00",x"3d"),
  3867 => (x"00",x"00",x"00",x"35"),
  3868 => (x"00",x"00",x"00",x"34"),
  3869 => (x"00",x"75",x"00",x"3e"),
  3870 => (x"00",x"00",x"00",x"32"),
  3871 => (x"00",x"00",x"00",x"33"),
  3872 => (x"00",x"6b",x"00",x"3c"),
  3873 => (x"00",x"00",x"00",x"2a"),
  3874 => (x"00",x"7d",x"00",x"46"),
  3875 => (x"00",x"73",x"00",x"43"),
  3876 => (x"00",x"69",x"00",x"3b"),
  3877 => (x"00",x"ca",x"00",x"45"),
  3878 => (x"00",x"70",x"00",x"3a"),
  3879 => (x"00",x"72",x"00",x"42"),
  3880 => (x"00",x"74",x"00",x"44"),
  3881 => (x"00",x"00",x"00",x"31"),
  3882 => (x"00",x"00",x"00",x"55"),
  3883 => (x"00",x"7c",x"00",x"4d"),
  3884 => (x"00",x"7a",x"00",x"4b"),
  3885 => (x"00",x"00",x"00",x"7b"),
  3886 => (x"00",x"71",x"00",x"49"),
  3887 => (x"00",x"84",x"00",x"4c"),
  3888 => (x"00",x"77",x"00",x"54"),
  3889 => (x"00",x"00",x"00",x"41"),
  3890 => (x"00",x"00",x"00",x"61"),
  3891 => (x"00",x"7c",x"00",x"5b"),
  3892 => (x"00",x"00",x"00",x"52"),
  3893 => (x"00",x"00",x"00",x"f1"),
  3894 => (x"00",x"00",x"02",x"59"),
  3895 => (x"00",x"5d",x"00",x"0e"),
  3896 => (x"00",x"00",x"00",x"5d"),
  3897 => (x"00",x"79",x"00",x"4a"),
  3898 => (x"00",x"00",x"00",x"16"),
  3899 => (x"00",x"07",x"00",x"76"),
  3900 => (x"00",x"0d",x"04",x"14"),
  3901 => (x"00",x"00",x"00",x"1e"),
  3902 => (x"00",x"00",x"00",x"29"),
  3903 => (x"00",x"00",x"00",x"11"),
  3904 => (x"00",x"00",x"00",x"15"),
  3905 => (x"00",x"00",x"40",x"00"),
  3906 => (x"00",x"00",x"3d",x"24"),
  3907 => (x"08",x"82",x"ff",x"01"),
  3908 => (x"64",x"f3",x"c8",x"f3"),
  3909 => (x"01",x"f2",x"50",x"f3"),
  3910 => (x"00",x"f4",x"01",x"81"),
  3911 => (x"00",x"00",x"3f",x"90"),
  3912 => (x"00",x"00",x"3f",x"9c"),
  3913 => (x"72",x"61",x"74",x"41"),
  3914 => (x"54",x"53",x"20",x"69"),
  3915 => (x"31",x"50",x"3b",x"3b"),
  3916 => (x"6f",x"74",x"53",x"2c"),
  3917 => (x"65",x"67",x"61",x"72"),
  3918 => (x"53",x"31",x"50",x"3b"),
  3919 => (x"53",x"2c",x"55",x"30"),
  3920 => (x"46",x"2c",x"20",x"54"),
  3921 => (x"70",x"70",x"6f",x"6c"),
  3922 => (x"3a",x"41",x"20",x"79"),
  3923 => (x"53",x"31",x"50",x"3b"),
  3924 => (x"53",x"2c",x"55",x"31"),
  3925 => (x"46",x"2c",x"20",x"54"),
  3926 => (x"70",x"70",x"6f",x"6c"),
  3927 => (x"3a",x"42",x"20",x"79"),
  3928 => (x"4f",x"31",x"50",x"3b"),
  3929 => (x"57",x"2c",x"37",x"36"),
  3930 => (x"65",x"74",x"69",x"72"),
  3931 => (x"6f",x"72",x"70",x"20"),
  3932 => (x"74",x"63",x"65",x"74"),
  3933 => (x"66",x"66",x"4f",x"2c"),
  3934 => (x"2c",x"3a",x"41",x"2c"),
  3935 => (x"42",x"2c",x"3a",x"42"),
  3936 => (x"3b",x"68",x"74",x"6f"),
  3937 => (x"41",x"4f",x"31",x"50"),
  3938 => (x"61",x"48",x"2c",x"42"),
  3939 => (x"64",x"20",x"64",x"72"),
  3940 => (x"73",x"6b",x"73",x"69"),
  3941 => (x"6e",x"6f",x"4e",x"2c"),
  3942 => (x"6e",x"55",x"2c",x"65"),
  3943 => (x"30",x"20",x"74",x"69"),
  3944 => (x"69",x"6e",x"55",x"2c"),
  3945 => (x"2c",x"31",x"20",x"74"),
  3946 => (x"68",x"74",x"6f",x"42"),
  3947 => (x"53",x"31",x"50",x"3b"),
  3948 => (x"48",x"2c",x"55",x"32"),
  3949 => (x"48",x"56",x"46",x"44"),
  3950 => (x"61",x"48",x"2c",x"44"),
  3951 => (x"69",x"66",x"64",x"72"),
  3952 => (x"30",x"20",x"65",x"6c"),
  3953 => (x"53",x"31",x"50",x"3b"),
  3954 => (x"48",x"2c",x"55",x"33"),
  3955 => (x"48",x"56",x"46",x"44"),
  3956 => (x"61",x"48",x"2c",x"44"),
  3957 => (x"69",x"66",x"64",x"72"),
  3958 => (x"31",x"20",x"65",x"6c"),
  3959 => (x"2c",x"32",x"50",x"3b"),
  3960 => (x"74",x"73",x"79",x"53"),
  3961 => (x"50",x"3b",x"6d",x"65"),
  3962 => (x"4f",x"4e",x"4f",x"32"),
  3963 => (x"69",x"68",x"43",x"2c"),
  3964 => (x"74",x"65",x"73",x"70"),
  3965 => (x"2c",x"54",x"53",x"2c"),
  3966 => (x"2c",x"45",x"54",x"53"),
  3967 => (x"61",x"67",x"65",x"4d"),
  3968 => (x"2c",x"45",x"54",x"53"),
  3969 => (x"72",x"45",x"54",x"53"),
  3970 => (x"73",x"64",x"69",x"6f"),
  3971 => (x"4f",x"32",x"50",x"3b"),
  3972 => (x"54",x"53",x"2c",x"4a"),
  3973 => (x"69",x"6c",x"42",x"20"),
  3974 => (x"72",x"65",x"74",x"74"),
  3975 => (x"66",x"66",x"4f",x"2c"),
  3976 => (x"3b",x"6e",x"4f",x"2c"),
  3977 => (x"31",x"4f",x"32",x"50"),
  3978 => (x"41",x"52",x"2c",x"33"),
  3979 => (x"6e",x"28",x"20",x"4d"),
  3980 => (x"20",x"64",x"65",x"65"),
  3981 => (x"64",x"72",x"61",x"48"),
  3982 => (x"73",x"65",x"52",x"20"),
  3983 => (x"2c",x"29",x"74",x"65"),
  3984 => (x"4b",x"32",x"31",x"35"),
  3985 => (x"42",x"4d",x"31",x"2c"),
  3986 => (x"42",x"4d",x"32",x"2c"),
  3987 => (x"42",x"4d",x"34",x"2c"),
  3988 => (x"42",x"4d",x"38",x"2c"),
  3989 => (x"4d",x"34",x"31",x"2c"),
  3990 => (x"32",x"50",x"3b",x"42"),
  3991 => (x"4d",x"49",x"2c",x"46"),
  3992 => (x"4d",x"4f",x"52",x"47"),
  3993 => (x"61",x"6f",x"4c",x"2c"),
  3994 => (x"4f",x"52",x"20",x"64"),
  3995 => (x"32",x"50",x"3b",x"4d"),
  3996 => (x"49",x"42",x"2c",x"46"),
  3997 => (x"43",x"54",x"53",x"4e"),
  3998 => (x"61",x"6f",x"4c",x"2c"),
  3999 => (x"61",x"43",x"20",x"64"),
  4000 => (x"69",x"72",x"74",x"72"),
  4001 => (x"3b",x"65",x"67",x"64"),
  4002 => (x"53",x"2c",x"33",x"50"),
  4003 => (x"64",x"6e",x"75",x"6f"),
  4004 => (x"56",x"20",x"26",x"20"),
  4005 => (x"6f",x"65",x"64",x"69"),
  4006 => (x"4f",x"33",x"50",x"3b"),
  4007 => (x"69",x"56",x"2c",x"38"),
  4008 => (x"20",x"6f",x"65",x"64"),
  4009 => (x"65",x"64",x"6f",x"6d"),
  4010 => (x"6e",x"6f",x"4d",x"2c"),
  4011 => (x"6f",x"43",x"2c",x"6f"),
  4012 => (x"72",x"75",x"6f",x"6c"),
  4013 => (x"4f",x"33",x"50",x"3b"),
  4014 => (x"69",x"56",x"2c",x"53"),
  4015 => (x"67",x"6e",x"69",x"6b"),
  4016 => (x"31",x"4d",x"53",x"2f"),
  4017 => (x"4f",x"2c",x"34",x"39"),
  4018 => (x"4f",x"2c",x"66",x"66"),
  4019 => (x"33",x"50",x"3b",x"6e"),
  4020 => (x"2c",x"4c",x"4b",x"4f"),
  4021 => (x"6e",x"61",x"63",x"53"),
  4022 => (x"65",x"6e",x"69",x"6c"),
  4023 => (x"66",x"4f",x"2c",x"73"),
  4024 => (x"35",x"32",x"2c",x"66"),
  4025 => (x"30",x"35",x"2c",x"25"),
  4026 => (x"35",x"37",x"2c",x"25"),
  4027 => (x"33",x"50",x"3b",x"25"),
  4028 => (x"43",x"2c",x"54",x"4f"),
  4029 => (x"6f",x"70",x"6d",x"6f"),
  4030 => (x"65",x"74",x"69",x"73"),
  4031 => (x"65",x"6c",x"62",x"20"),
  4032 => (x"4f",x"2c",x"64",x"6e"),
  4033 => (x"4f",x"2c",x"66",x"66"),
  4034 => (x"33",x"50",x"3b",x"6e"),
  4035 => (x"53",x"2c",x"4d",x"4f"),
  4036 => (x"65",x"72",x"65",x"74"),
  4037 => (x"6f",x"73",x"20",x"6f"),
  4038 => (x"2c",x"64",x"6e",x"75"),
  4039 => (x"2c",x"66",x"66",x"4f"),
  4040 => (x"50",x"3b",x"6e",x"4f"),
  4041 => (x"2c",x"55",x"4f",x"33"),
  4042 => (x"69",x"65",x"74",x"53"),
  4043 => (x"72",x"65",x"62",x"6e"),
  4044 => (x"6f",x"64",x"20",x"67"),
  4045 => (x"65",x"6c",x"67",x"6e"),
  4046 => (x"66",x"66",x"4f",x"2c"),
  4047 => (x"3b",x"6e",x"4f",x"2c"),
  4048 => (x"43",x"2c",x"43",x"53"),
  4049 => (x"4c",x"2c",x"47",x"46"),
  4050 => (x"20",x"64",x"61",x"6f"),
  4051 => (x"66",x"6e",x"6f",x"63"),
  4052 => (x"53",x"3b",x"67",x"69"),
  4053 => (x"46",x"43",x"2c",x"44"),
  4054 => (x"61",x"53",x"2c",x"47"),
  4055 => (x"63",x"20",x"65",x"76"),
  4056 => (x"69",x"66",x"6e",x"6f"),
  4057 => (x"30",x"54",x"3b",x"67"),
  4058 => (x"73",x"65",x"52",x"2c"),
  4059 => (x"28",x"20",x"74",x"65"),
  4060 => (x"64",x"6c",x"6f",x"48"),
  4061 => (x"72",x"6f",x"66",x"20"),
  4062 => (x"72",x"61",x"68",x"20"),
  4063 => (x"65",x"72",x"20",x"64"),
  4064 => (x"29",x"74",x"65",x"73"),
  4065 => (x"76",x"2c",x"56",x"3b"),
  4066 => (x"30",x"34",x"2e",x"33"),
  4067 => (x"00",x"00",x"00",x"2e"),
  4068 => (x"20",x"53",x"4f",x"54"),
  4069 => (x"20",x"20",x"20",x"20"),
  4070 => (x"00",x"47",x"4d",x"49"),
  4071 => (x"54",x"53",x"49",x"4d"),
  4072 => (x"20",x"59",x"52",x"45"),
  4073 => (x"00",x"47",x"46",x"43"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

