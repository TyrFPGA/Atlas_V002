library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dcfac287",
    12 => x"86c0c54e",
    13 => x"49dcfac2",
    14 => x"48e8e7c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087eae3",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfe8e7",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"e7c21e73",
   183 => x"78c148e8",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"ece7c287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58f0e7c2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49f0e7c2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97f0e7",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97f7e7",
   291 => x"c231d049",
   292 => x"bf97f8e7",
   293 => x"7232c84a",
   294 => x"f9e7c2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"e7c287e7",
   300 => x"49bf97f9",
   301 => x"99c631c1",
   302 => x"97fae7c2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97f5e7",
   306 => x"9dcf4d4a",
   307 => x"97f6e7c2",
   308 => x"9ac34abf",
   309 => x"e7c232ca",
   310 => x"4bbf97f7",
   311 => x"b27333c2",
   312 => x"97f8e7c2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"f0c286f8",
   329 => x"78c048d6",
   330 => x"1ecee8c2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"ddf2c07e",
   337 => x"e9c249bf",
   338 => x"c8714ac4",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfd9f2",
   343 => x"4ae0e9c2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"efc287fd",
   349 => x"c24dbfd4",
   350 => x"bf9fccf0",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"d4efc287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"e8c287e3",
   359 => x"49751ece",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfd9f2",
   365 => x"4ae0e9c2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148d6f0",
   370 => x"c087da78",
   371 => x"49bfddf2",
   372 => x"4ac4e9c2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"ccf0c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"f0c287cd",
   381 => x"49bf97cd",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97cee8c2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97d9e8c2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97dae8",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97dbe8c2",
   400 => x"f0c248bf",
   401 => x"4c7058d2",
   402 => x"c288c148",
   403 => x"c258d6f0",
   404 => x"bf97dce8",
   405 => x"c2817549",
   406 => x"bf97dde8",
   407 => x"7232c84a",
   408 => x"f4c27ea1",
   409 => x"786e48e3",
   410 => x"97dee8c2",
   411 => x"a6c848bf",
   412 => x"d6f0c258",
   413 => x"cfc202bf",
   414 => x"d9f2c087",
   415 => x"e9c249bf",
   416 => x"c8714ae0",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbfcef0",
   422 => x"5cf7f4c2",
   423 => x"97f3e8c2",
   424 => x"31c849bf",
   425 => x"97f2e8c2",
   426 => x"49a14abf",
   427 => x"97f4e8c2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97f5e8",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"e3f4c291",
   434 => x"f4c281bf",
   435 => x"e8c259eb",
   436 => x"4abf97fb",
   437 => x"e8c232c8",
   438 => x"4bbf97fa",
   439 => x"e8c24aa2",
   440 => x"4bbf97fc",
   441 => x"a27333d0",
   442 => x"fde8c24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"f4c24aa2",
   446 => x"8ac25aef",
   447 => x"f4c29274",
   448 => x"a17248ef",
   449 => x"87c1c178",
   450 => x"97e0e8c2",
   451 => x"31c849bf",
   452 => x"97dfe8c2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259f7f4",
   457 => x"bf97e5e8",
   458 => x"c232c84a",
   459 => x"bf97e4e8",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5af3f4c2",
   463 => x"48ebf4c2",
   464 => x"f4c278c0",
   465 => x"a17248e7",
   466 => x"f7f4c278",
   467 => x"ebf4c248",
   468 => x"f4c278bf",
   469 => x"f4c248fb",
   470 => x"c278bfef",
   471 => x"02bfd6f0",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bff3f4c2",
   476 => x"7030c448",
   477 => x"daf0c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfd6f0",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"f4c29dff",
   491 => x"c083bfe3",
   492 => x"abbfd5f2",
   493 => x"c087d902",
   494 => x"c25bd9f2",
   495 => x"731ecee8",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfd6f0c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981cee8",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"cee8c291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c0c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087e9c2",
   521 => x"4949c11e",
   522 => x"c487d3ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4adef0c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d1c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cec102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfd6f0",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"486e7ec0",
   556 => x"80bf66c4",
   557 => x"780866c4",
   558 => x"a4cc7cc0",
   559 => x"bf66c449",
   560 => x"49a4d079",
   561 => x"48c179c0",
   562 => x"48c087c2",
   563 => x"eefa8ef8",
   564 => x"5b5e0e87",
   565 => x"4c710e5c",
   566 => x"cbc1029c",
   567 => x"49a4c887",
   568 => x"c3c10269",
   569 => x"cc496c87",
   570 => x"80714866",
   571 => x"7058a6d0",
   572 => x"d2f0c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e5c002",
   576 => x"6b4ba4c4",
   577 => x"87fff949",
   578 => x"f0c27b70",
   579 => x"6c49bfce",
   580 => x"cc7c7181",
   581 => x"f0c2b966",
   582 => x"ff4abfd2",
   583 => x"719972ba",
   584 => x"dbff0599",
   585 => x"7c66cc87",
   586 => x"1e87d6f9",
   587 => x"4b711e73",
   588 => x"87c7029b",
   589 => x"6949a3c8",
   590 => x"c087c505",
   591 => x"87f6c048",
   592 => x"bfe7f4c2",
   593 => x"4aa3c449",
   594 => x"8ac24a6a",
   595 => x"bfcef0c2",
   596 => x"49a17292",
   597 => x"bfd2f0c2",
   598 => x"729a6b4a",
   599 => x"f2c049a1",
   600 => x"66c859d9",
   601 => x"e6ea711e",
   602 => x"7086c487",
   603 => x"87c40598",
   604 => x"87c248c0",
   605 => x"caf848c1",
   606 => x"1e731e87",
   607 => x"029b4b71",
   608 => x"a3c887c7",
   609 => x"c5056949",
   610 => x"c048c087",
   611 => x"f4c287f6",
   612 => x"c449bfe7",
   613 => x"4a6a4aa3",
   614 => x"f0c28ac2",
   615 => x"7292bfce",
   616 => x"f0c249a1",
   617 => x"6b4abfd2",
   618 => x"49a1729a",
   619 => x"59d9f2c0",
   620 => x"711e66c8",
   621 => x"c487d1e6",
   622 => x"05987086",
   623 => x"48c087c4",
   624 => x"48c187c2",
   625 => x"0e87fcf6",
   626 => x"5d5c5b5e",
   627 => x"4b711e0e",
   628 => x"734d66d4",
   629 => x"ccc1029b",
   630 => x"49a3c887",
   631 => x"c4c10269",
   632 => x"4ca3d087",
   633 => x"bfd2f0c2",
   634 => x"6cb9ff49",
   635 => x"d47e994a",
   636 => x"cd06a966",
   637 => x"7c7bc087",
   638 => x"c44aa3cc",
   639 => x"796a49a3",
   640 => x"497287ca",
   641 => x"d499c0f8",
   642 => x"8d714d66",
   643 => x"29c94975",
   644 => x"49731e71",
   645 => x"c287fafa",
   646 => x"731ecee8",
   647 => x"87cbfc49",
   648 => x"66d486c8",
   649 => x"d6f5267c",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"c287e4c0",
   653 => x"735bfbf4",
   654 => x"c28ac24a",
   655 => x"49bfcef0",
   656 => x"e7f4c292",
   657 => x"807248bf",
   658 => x"58fff4c2",
   659 => x"30c44871",
   660 => x"58def0c2",
   661 => x"c287edc0",
   662 => x"c248f7f4",
   663 => x"78bfebf4",
   664 => x"48fbf4c2",
   665 => x"bfeff4c2",
   666 => x"d6f0c278",
   667 => x"87c902bf",
   668 => x"bfcef0c2",
   669 => x"c731c449",
   670 => x"f3f4c287",
   671 => x"31c449bf",
   672 => x"59def0c2",
   673 => x"0e87fcf3",
   674 => x"0e5c5b5e",
   675 => x"4bc04a71",
   676 => x"c0029a72",
   677 => x"a2da87e0",
   678 => x"4b699f49",
   679 => x"bfd6f0c2",
   680 => x"d487cf02",
   681 => x"699f49a2",
   682 => x"ffc04c49",
   683 => x"34d09cff",
   684 => x"4cc087c2",
   685 => x"4973b374",
   686 => x"f387eefd",
   687 => x"5e0e87c3",
   688 => x"0e5d5c5b",
   689 => x"4a7186f4",
   690 => x"9a727ec0",
   691 => x"c287d802",
   692 => x"c048cae8",
   693 => x"c2e8c278",
   694 => x"fbf4c248",
   695 => x"e8c278bf",
   696 => x"f4c248c6",
   697 => x"c278bff7",
   698 => x"c048ebf0",
   699 => x"daf0c250",
   700 => x"e8c249bf",
   701 => x"714abfca",
   702 => x"c9c403aa",
   703 => x"cf497287",
   704 => x"e9c00599",
   705 => x"d5f2c087",
   706 => x"c2e8c248",
   707 => x"e8c278bf",
   708 => x"e8c21ece",
   709 => x"c249bfc2",
   710 => x"c148c2e8",
   711 => x"e37178a1",
   712 => x"86c487ed",
   713 => x"48d1f2c0",
   714 => x"78cee8c2",
   715 => x"f2c087cc",
   716 => x"c048bfd1",
   717 => x"f2c080e0",
   718 => x"e8c258d5",
   719 => x"c148bfca",
   720 => x"cee8c280",
   721 => x"0c912758",
   722 => x"97bf0000",
   723 => x"029d4dbf",
   724 => x"c387e3c2",
   725 => x"c202ade5",
   726 => x"f2c087dc",
   727 => x"cb4bbfd1",
   728 => x"4c1149a3",
   729 => x"c105accf",
   730 => x"497587d2",
   731 => x"89c199df",
   732 => x"f0c291cd",
   733 => x"a3c181de",
   734 => x"c351124a",
   735 => x"51124aa3",
   736 => x"124aa3c5",
   737 => x"4aa3c751",
   738 => x"a3c95112",
   739 => x"ce51124a",
   740 => x"51124aa3",
   741 => x"124aa3d0",
   742 => x"4aa3d251",
   743 => x"a3d45112",
   744 => x"d651124a",
   745 => x"51124aa3",
   746 => x"124aa3d8",
   747 => x"4aa3dc51",
   748 => x"a3de5112",
   749 => x"c151124a",
   750 => x"87fac07e",
   751 => x"99c84974",
   752 => x"87ebc005",
   753 => x"99d04974",
   754 => x"dc87d105",
   755 => x"cbc00266",
   756 => x"dc497387",
   757 => x"98700f66",
   758 => x"87d3c002",
   759 => x"c6c0056e",
   760 => x"def0c287",
   761 => x"c050c048",
   762 => x"48bfd1f2",
   763 => x"c287ddc2",
   764 => x"c048ebf0",
   765 => x"f0c27e50",
   766 => x"c249bfda",
   767 => x"4abfcae8",
   768 => x"fb04aa71",
   769 => x"f4c287f7",
   770 => x"c005bffb",
   771 => x"f0c287c8",
   772 => x"c102bfd6",
   773 => x"e8c287f4",
   774 => x"ed49bfc6",
   775 => x"e8c287e9",
   776 => x"a6c458ca",
   777 => x"c6e8c248",
   778 => x"f0c278bf",
   779 => x"c002bfd6",
   780 => x"66c487d8",
   781 => x"ffffcf49",
   782 => x"a999f8ff",
   783 => x"87c5c002",
   784 => x"e1c04cc0",
   785 => x"c04cc187",
   786 => x"66c487dc",
   787 => x"f8ffcf49",
   788 => x"c002a999",
   789 => x"a6c887c8",
   790 => x"c078c048",
   791 => x"a6c887c5",
   792 => x"c878c148",
   793 => x"9c744c66",
   794 => x"87dec005",
   795 => x"c24966c4",
   796 => x"cef0c289",
   797 => x"f4c291bf",
   798 => x"7148bfe7",
   799 => x"c6e8c280",
   800 => x"cae8c258",
   801 => x"f978c048",
   802 => x"48c087e3",
   803 => x"eeeb8ef4",
   804 => x"00000087",
   805 => x"ffffff00",
   806 => x"000ca1ff",
   807 => x"000caa00",
   808 => x"54414600",
   809 => x"20203233",
   810 => x"41460020",
   811 => x"20363154",
   812 => x"1e002020",
   813 => x"c348d4ff",
   814 => x"486878ff",
   815 => x"ff1e4f26",
   816 => x"ffc348d4",
   817 => x"48d0ff78",
   818 => x"ff78e1c0",
   819 => x"78d448d4",
   820 => x"48fff4c2",
   821 => x"50bfd4ff",
   822 => x"ff1e4f26",
   823 => x"e0c048d0",
   824 => x"1e4f2678",
   825 => x"7087ccff",
   826 => x"c6029949",
   827 => x"a9fbc087",
   828 => x"7187f105",
   829 => x"0e4f2648",
   830 => x"0e5c5b5e",
   831 => x"4cc04b71",
   832 => x"7087f0fe",
   833 => x"c0029949",
   834 => x"ecc087f9",
   835 => x"f2c002a9",
   836 => x"a9fbc087",
   837 => x"87ebc002",
   838 => x"acb766cc",
   839 => x"d087c703",
   840 => x"87c20266",
   841 => x"99715371",
   842 => x"c187c202",
   843 => x"87c3fe84",
   844 => x"02994970",
   845 => x"ecc087cd",
   846 => x"87c702a9",
   847 => x"05a9fbc0",
   848 => x"d087d5ff",
   849 => x"87c30266",
   850 => x"c07b97c0",
   851 => x"c405a9ec",
   852 => x"c54a7487",
   853 => x"c04a7487",
   854 => x"48728a0a",
   855 => x"4d2687c2",
   856 => x"4b264c26",
   857 => x"fd1e4f26",
   858 => x"497087c9",
   859 => x"aaf0c04a",
   860 => x"c087c904",
   861 => x"c301aaf9",
   862 => x"8af0c087",
   863 => x"04aac1c1",
   864 => x"dac187c9",
   865 => x"87c301aa",
   866 => x"728af7c0",
   867 => x"0e4f2648",
   868 => x"5d5c5b5e",
   869 => x"7186f80e",
   870 => x"c04dc04b",
   871 => x"bf97e8f9",
   872 => x"05a9df49",
   873 => x"c887eec0",
   874 => x"699749a3",
   875 => x"a9c3c149",
   876 => x"c987dd05",
   877 => x"699749a3",
   878 => x"a9c6c149",
   879 => x"ca87d105",
   880 => x"699749a3",
   881 => x"a9c7c149",
   882 => x"c187c505",
   883 => x"87d3c248",
   884 => x"cec248c0",
   885 => x"87e6fb87",
   886 => x"f9c04cc0",
   887 => x"49bf97e8",
   888 => x"cf04a9c0",
   889 => x"87fbfb87",
   890 => x"f9c084c1",
   891 => x"49bf97e8",
   892 => x"87f106ac",
   893 => x"97e8f9c0",
   894 => x"87cf02bf",
   895 => x"7087f4fa",
   896 => x"c6029949",
   897 => x"a9ecc087",
   898 => x"c087f105",
   899 => x"87e3fa4c",
   900 => x"defa7e70",
   901 => x"58a6c887",
   902 => x"7087d8fa",
   903 => x"c884c14a",
   904 => x"699749a3",
   905 => x"05a96e49",
   906 => x"a3c987da",
   907 => x"49699749",
   908 => x"05a966c4",
   909 => x"a3ca87ce",
   910 => x"49699749",
   911 => x"87c405aa",
   912 => x"87d44dc1",
   913 => x"ecc0486e",
   914 => x"87c802a8",
   915 => x"fbc0486e",
   916 => x"87c405a8",
   917 => x"4dc14cc0",
   918 => x"fe029d75",
   919 => x"f9f987ef",
   920 => x"f8487487",
   921 => x"87f6fb8e",
   922 => x"5b5e0e00",
   923 => x"f80e5d5c",
   924 => x"ff7e7186",
   925 => x"1e6e4bd4",
   926 => x"49c4f5c2",
   927 => x"c487fae5",
   928 => x"02987086",
   929 => x"c187eac4",
   930 => x"4dbfcee7",
   931 => x"fefb496e",
   932 => x"58a6c887",
   933 => x"c5059870",
   934 => x"48a6c487",
   935 => x"d0ff78c1",
   936 => x"c178c548",
   937 => x"66c47bd5",
   938 => x"c689c149",
   939 => x"cce7c131",
   940 => x"484abf97",
   941 => x"7b70b071",
   942 => x"c448d0ff",
   943 => x"fff4c278",
   944 => x"d049bf97",
   945 => x"87d70299",
   946 => x"d6c178c5",
   947 => x"c34ac07b",
   948 => x"82c17bff",
   949 => x"04aae0c0",
   950 => x"d0ff87f5",
   951 => x"c378c448",
   952 => x"d0ff7bff",
   953 => x"c178c548",
   954 => x"7bc17bd3",
   955 => x"b7c078c4",
   956 => x"ebc206ad",
   957 => x"ccf5c287",
   958 => x"9c8d4cbf",
   959 => x"87c2c202",
   960 => x"7ecee8c2",
   961 => x"c848a6c4",
   962 => x"c08c78c0",
   963 => x"c603acb7",
   964 => x"a4c0c887",
   965 => x"c24cc078",
   966 => x"bf97fff4",
   967 => x"0299d049",
   968 => x"1ec087d0",
   969 => x"49c4f5c2",
   970 => x"c487c0e8",
   971 => x"c04a7086",
   972 => x"e8c287f5",
   973 => x"f5c21ece",
   974 => x"eee749c4",
   975 => x"7086c487",
   976 => x"48d0ff4a",
   977 => x"c178c5c8",
   978 => x"976e7bd4",
   979 => x"486e7bbf",
   980 => x"7e7080c1",
   981 => x"c14866c4",
   982 => x"58a6c888",
   983 => x"ff059870",
   984 => x"d0ff87e8",
   985 => x"7278c448",
   986 => x"87c5059a",
   987 => x"c2c148c0",
   988 => x"c21ec187",
   989 => x"e549c4f5",
   990 => x"86c487d7",
   991 => x"fd059c74",
   992 => x"b7c087fe",
   993 => x"87d106ad",
   994 => x"48c4f5c2",
   995 => x"80d078c0",
   996 => x"80f478c0",
   997 => x"bfd0f5c2",
   998 => x"adb7c078",
   999 => x"87d5fd01",
  1000 => x"c548d0ff",
  1001 => x"7bd3c178",
  1002 => x"78c47bc0",
  1003 => x"c2c048c1",
  1004 => x"f848c087",
  1005 => x"264d268e",
  1006 => x"264b264c",
  1007 => x"5b5e0e4f",
  1008 => x"1e0e5d5c",
  1009 => x"4cc04b71",
  1010 => x"c004ab4d",
  1011 => x"f6c087e8",
  1012 => x"9d751ecf",
  1013 => x"c087c402",
  1014 => x"c187c24a",
  1015 => x"eb49724a",
  1016 => x"86c487dc",
  1017 => x"84c17e70",
  1018 => x"87c2056e",
  1019 => x"85c14c73",
  1020 => x"ff06ac73",
  1021 => x"486e87d8",
  1022 => x"87f9fe26",
  1023 => x"5c5b5e0e",
  1024 => x"cc4b710e",
  1025 => x"e8c00266",
  1026 => x"f0c04c87",
  1027 => x"e8c0028c",
  1028 => x"c14a7487",
  1029 => x"e0c0028a",
  1030 => x"dc028a87",
  1031 => x"d8028a87",
  1032 => x"8ae0c087",
  1033 => x"87e5c002",
  1034 => x"c0028ac1",
  1035 => x"eac087e7",
  1036 => x"f8497387",
  1037 => x"e2c087f3",
  1038 => x"c01e7487",
  1039 => x"cedec149",
  1040 => x"731e7487",
  1041 => x"c6dec149",
  1042 => x"ce86c887",
  1043 => x"c1497387",
  1044 => x"c687ebe0",
  1045 => x"c1497387",
  1046 => x"fd87dde1",
  1047 => x"5e0e87d9",
  1048 => x"0e5d5c5b",
  1049 => x"494c711e",
  1050 => x"f5c291de",
  1051 => x"85714dec",
  1052 => x"c1026d97",
  1053 => x"f5c287dd",
  1054 => x"7449bfd8",
  1055 => x"fcfc7181",
  1056 => x"487e7087",
  1057 => x"f2c00298",
  1058 => x"e0f5c287",
  1059 => x"cb4a704b",
  1060 => x"d2c0ff49",
  1061 => x"cb4b7487",
  1062 => x"c3e8c193",
  1063 => x"c183c483",
  1064 => x"747bd7c3",
  1065 => x"fec2c149",
  1066 => x"c17b7587",
  1067 => x"bf97cde7",
  1068 => x"f5c21e49",
  1069 => x"c3fd49e0",
  1070 => x"7486c487",
  1071 => x"e6c2c149",
  1072 => x"c149c087",
  1073 => x"c287c5c4",
  1074 => x"c048c0f5",
  1075 => x"c049c178",
  1076 => x"2687e5e0",
  1077 => x"4c87defb",
  1078 => x"6964616f",
  1079 => x"2e2e676e",
  1080 => x"731e002e",
  1081 => x"494a711e",
  1082 => x"bfd8f5c2",
  1083 => x"ccfb7181",
  1084 => x"9b4b7087",
  1085 => x"4987c402",
  1086 => x"c287cce6",
  1087 => x"c048d8f5",
  1088 => x"df49c178",
  1089 => x"f0fa87f2",
  1090 => x"49c01e87",
  1091 => x"87fcc2c1",
  1092 => x"711e4f26",
  1093 => x"91cb494a",
  1094 => x"81c3e8c1",
  1095 => x"481181c8",
  1096 => x"58c4f5c2",
  1097 => x"48d8f5c2",
  1098 => x"49c178c0",
  1099 => x"2687c9df",
  1100 => x"99711e4f",
  1101 => x"c187d202",
  1102 => x"c048d8e9",
  1103 => x"c180f750",
  1104 => x"c140d2c4",
  1105 => x"ce78f1e7",
  1106 => x"d4e9c187",
  1107 => x"d2e7c148",
  1108 => x"c180fc78",
  1109 => x"2678c9c4",
  1110 => x"5b5e0e4f",
  1111 => x"f40e5d5c",
  1112 => x"cee8c286",
  1113 => x"c44cc04d",
  1114 => x"78c048a6",
  1115 => x"bfd8f5c2",
  1116 => x"06a8c048",
  1117 => x"c287c0c1",
  1118 => x"9848cee8",
  1119 => x"87f7c002",
  1120 => x"1ecff6c0",
  1121 => x"c70266c8",
  1122 => x"48a6c487",
  1123 => x"87c578c0",
  1124 => x"c148a6c4",
  1125 => x"4966c478",
  1126 => x"c487e3e4",
  1127 => x"c14d7086",
  1128 => x"4866c484",
  1129 => x"a6c880c1",
  1130 => x"d8f5c258",
  1131 => x"c603acbf",
  1132 => x"059d7587",
  1133 => x"c087c9ff",
  1134 => x"029d754c",
  1135 => x"c087dcc3",
  1136 => x"c81ecff6",
  1137 => x"87c70266",
  1138 => x"c048a6cc",
  1139 => x"cc87c578",
  1140 => x"78c148a6",
  1141 => x"e34966cc",
  1142 => x"86c487e4",
  1143 => x"98487e70",
  1144 => x"87e4c202",
  1145 => x"9781cb49",
  1146 => x"99d04969",
  1147 => x"87d4c102",
  1148 => x"91cb4974",
  1149 => x"81c3e8c1",
  1150 => x"79e2c3c1",
  1151 => x"ffc381c8",
  1152 => x"de497451",
  1153 => x"ecf5c291",
  1154 => x"c285714d",
  1155 => x"c17d97c1",
  1156 => x"e0c049a5",
  1157 => x"def0c251",
  1158 => x"d202bf97",
  1159 => x"c284c187",
  1160 => x"f0c24ba5",
  1161 => x"49db4ade",
  1162 => x"87fbf9fe",
  1163 => x"cd87d9c1",
  1164 => x"51c049a5",
  1165 => x"a5c284c1",
  1166 => x"cb4a6e4b",
  1167 => x"e6f9fe49",
  1168 => x"87c4c187",
  1169 => x"91cb4974",
  1170 => x"81c3e8c1",
  1171 => x"79dec1c1",
  1172 => x"97def0c2",
  1173 => x"87d802bf",
  1174 => x"91de4974",
  1175 => x"f5c284c1",
  1176 => x"83714bec",
  1177 => x"4adef0c2",
  1178 => x"f8fe49dd",
  1179 => x"87d887f9",
  1180 => x"93de4b74",
  1181 => x"83ecf5c2",
  1182 => x"c049a3cb",
  1183 => x"7384c151",
  1184 => x"49cb4a6e",
  1185 => x"87dff8fe",
  1186 => x"c14866c4",
  1187 => x"58a6c880",
  1188 => x"c003acc7",
  1189 => x"056e87c5",
  1190 => x"7487e4fc",
  1191 => x"f48ef448",
  1192 => x"731e87d3",
  1193 => x"494b711e",
  1194 => x"e8c191cb",
  1195 => x"a1c881c3",
  1196 => x"cce7c14a",
  1197 => x"c9501248",
  1198 => x"f9c04aa1",
  1199 => x"501248e8",
  1200 => x"e7c181ca",
  1201 => x"501148cd",
  1202 => x"97cde7c1",
  1203 => x"c01e49bf",
  1204 => x"87e8f449",
  1205 => x"48c0f5c2",
  1206 => x"49c178de",
  1207 => x"2687d9d8",
  1208 => x"0e87d6f3",
  1209 => x"5d5c5b5e",
  1210 => x"7186f40e",
  1211 => x"91cb494d",
  1212 => x"81c3e8c1",
  1213 => x"ca4aa1c8",
  1214 => x"a6c47ea1",
  1215 => x"c8f9c248",
  1216 => x"976e78bf",
  1217 => x"66c44bbf",
  1218 => x"122c734c",
  1219 => x"58a6cc48",
  1220 => x"84c19c70",
  1221 => x"699781c9",
  1222 => x"04acb749",
  1223 => x"4cc087c2",
  1224 => x"4abf976e",
  1225 => x"724966c8",
  1226 => x"c4b9ff31",
  1227 => x"48749966",
  1228 => x"4a703072",
  1229 => x"c2b07148",
  1230 => x"c058ccf9",
  1231 => x"c087e8e6",
  1232 => x"87f4d649",
  1233 => x"f8c04975",
  1234 => x"8ef487dd",
  1235 => x"1e87e6f1",
  1236 => x"4b711e73",
  1237 => x"87cbfe49",
  1238 => x"c6fe4973",
  1239 => x"87d9f187",
  1240 => x"711e731e",
  1241 => x"4aa3c64b",
  1242 => x"87e3c002",
  1243 => x"d6028ac1",
  1244 => x"c1028a87",
  1245 => x"028a87e8",
  1246 => x"8a87cac1",
  1247 => x"87efc002",
  1248 => x"87d9028a",
  1249 => x"c787e9c1",
  1250 => x"87c6f649",
  1251 => x"c287ecc1",
  1252 => x"df48c0f5",
  1253 => x"d549c178",
  1254 => x"dec187de",
  1255 => x"d8f5c287",
  1256 => x"cbc102bf",
  1257 => x"88c14887",
  1258 => x"58dcf5c2",
  1259 => x"c287c1c1",
  1260 => x"02bfdcf5",
  1261 => x"c287f9c0",
  1262 => x"48bfd8f5",
  1263 => x"f5c280c1",
  1264 => x"ebc058dc",
  1265 => x"d8f5c287",
  1266 => x"89c649bf",
  1267 => x"59dcf5c2",
  1268 => x"03a9b7c0",
  1269 => x"f5c287da",
  1270 => x"78c048d8",
  1271 => x"f5c287d2",
  1272 => x"cb02bfdc",
  1273 => x"d8f5c287",
  1274 => x"80c648bf",
  1275 => x"58dcf5c2",
  1276 => x"c3d449c0",
  1277 => x"c0497387",
  1278 => x"ee87ecf5",
  1279 => x"5e0e87fb",
  1280 => x"0e5d5c5b",
  1281 => x"dc86d4ff",
  1282 => x"a6c859a6",
  1283 => x"c478c048",
  1284 => x"66c0c180",
  1285 => x"c180c478",
  1286 => x"c180c478",
  1287 => x"dcf5c278",
  1288 => x"c278c148",
  1289 => x"7ebfc0f5",
  1290 => x"a8de486e",
  1291 => x"f487c905",
  1292 => x"a6cc87e7",
  1293 => x"87dfd158",
  1294 => x"a8df486e",
  1295 => x"87eac105",
  1296 => x"4966fcc0",
  1297 => x"7e6981c4",
  1298 => x"48cce3c1",
  1299 => x"a1d0496e",
  1300 => x"7141204a",
  1301 => x"87f905aa",
  1302 => x"4866fcc0",
  1303 => x"78e2cac1",
  1304 => x"4966fcc0",
  1305 => x"51df81c9",
  1306 => x"4966fcc0",
  1307 => x"d3c181ca",
  1308 => x"66fcc051",
  1309 => x"c481cb49",
  1310 => x"a6c44aa1",
  1311 => x"71786a48",
  1312 => x"dce3c11e",
  1313 => x"4966c848",
  1314 => x"204aa1d0",
  1315 => x"05aa7141",
  1316 => x"492687f9",
  1317 => x"79e2cac1",
  1318 => x"df4aa1c9",
  1319 => x"c181ca52",
  1320 => x"a6c851d4",
  1321 => x"cf78c248",
  1322 => x"d1e087ed",
  1323 => x"87f3e087",
  1324 => x"7087c0e0",
  1325 => x"acfbc04c",
  1326 => x"87fdc102",
  1327 => x"c10566d8",
  1328 => x"fcc087ee",
  1329 => x"82c44a66",
  1330 => x"1e727e6a",
  1331 => x"48ece3c1",
  1332 => x"c84966c4",
  1333 => x"41204aa1",
  1334 => x"f905aa71",
  1335 => x"26511087",
  1336 => x"66fcc04a",
  1337 => x"e2cac148",
  1338 => x"c7496a78",
  1339 => x"c0517481",
  1340 => x"c84966fc",
  1341 => x"c051c181",
  1342 => x"c94966fc",
  1343 => x"c051c081",
  1344 => x"ca4966fc",
  1345 => x"c151c081",
  1346 => x"6a1ed81e",
  1347 => x"ff81c849",
  1348 => x"c887e4df",
  1349 => x"66c0c186",
  1350 => x"01a8c048",
  1351 => x"a6c887c7",
  1352 => x"cf78c148",
  1353 => x"66c0c187",
  1354 => x"d088c148",
  1355 => x"87c458a6",
  1356 => x"87efdeff",
  1357 => x"c248a6d0",
  1358 => x"029c7478",
  1359 => x"c887d4cd",
  1360 => x"c4c14866",
  1361 => x"cd03a866",
  1362 => x"a6dc87c9",
  1363 => x"e878c048",
  1364 => x"ff78c080",
  1365 => x"7087dcdd",
  1366 => x"acd0c14c",
  1367 => x"87d9c205",
  1368 => x"e07e66c4",
  1369 => x"a6c887c0",
  1370 => x"c6ddff58",
  1371 => x"c04c7087",
  1372 => x"c105acec",
  1373 => x"66c887ed",
  1374 => x"c091cb49",
  1375 => x"c48166fc",
  1376 => x"4d6a4aa1",
  1377 => x"c44aa1c8",
  1378 => x"c4c15266",
  1379 => x"dcff79d2",
  1380 => x"4c7087e1",
  1381 => x"87d9029c",
  1382 => x"02acfbc0",
  1383 => x"557487d3",
  1384 => x"87cfdcff",
  1385 => x"029c4c70",
  1386 => x"fbc087c7",
  1387 => x"edff05ac",
  1388 => x"55e0c087",
  1389 => x"c055c1c2",
  1390 => x"66d87d97",
  1391 => x"05a86e48",
  1392 => x"66c887db",
  1393 => x"a866cc48",
  1394 => x"c887ca04",
  1395 => x"80c14866",
  1396 => x"c858a6cc",
  1397 => x"4866cc87",
  1398 => x"a6d088c1",
  1399 => x"d2dbff58",
  1400 => x"c14c7087",
  1401 => x"c005acd0",
  1402 => x"66d487c8",
  1403 => x"d880c148",
  1404 => x"d0c158a6",
  1405 => x"e7fd02ac",
  1406 => x"4866c487",
  1407 => x"05a866d8",
  1408 => x"c087e2c9",
  1409 => x"c048a6e0",
  1410 => x"c0487478",
  1411 => x"7e7088fb",
  1412 => x"c9029848",
  1413 => x"cb4887e4",
  1414 => x"487e7088",
  1415 => x"cfc10298",
  1416 => x"88c94887",
  1417 => x"98487e70",
  1418 => x"87c0c402",
  1419 => x"7088c448",
  1420 => x"0298487e",
  1421 => x"4887cec0",
  1422 => x"7e7088c1",
  1423 => x"c3029848",
  1424 => x"d7c887ea",
  1425 => x"48a6dc87",
  1426 => x"ff78f0c0",
  1427 => x"7087e4d9",
  1428 => x"acecc04c",
  1429 => x"87c4c002",
  1430 => x"5ca6e0c0",
  1431 => x"02acecc0",
  1432 => x"ff87cdc0",
  1433 => x"7087ccd9",
  1434 => x"acecc04c",
  1435 => x"87f3ff05",
  1436 => x"02acecc0",
  1437 => x"ff87c4c0",
  1438 => x"c087f8d8",
  1439 => x"d01eca1e",
  1440 => x"91cb4966",
  1441 => x"4866c4c1",
  1442 => x"a6cc8071",
  1443 => x"4866c858",
  1444 => x"a6d080c4",
  1445 => x"bf66cc58",
  1446 => x"dad9ff49",
  1447 => x"de1ec187",
  1448 => x"bf66d41e",
  1449 => x"ced9ff49",
  1450 => x"7086d087",
  1451 => x"08c04849",
  1452 => x"a6e8c088",
  1453 => x"06a8c058",
  1454 => x"c087eec0",
  1455 => x"dd4866e4",
  1456 => x"e4c003a8",
  1457 => x"bf66c487",
  1458 => x"66e4c049",
  1459 => x"51e0c081",
  1460 => x"4966e4c0",
  1461 => x"66c481c1",
  1462 => x"c1c281bf",
  1463 => x"66e4c051",
  1464 => x"c481c249",
  1465 => x"c081bf66",
  1466 => x"c1486e51",
  1467 => x"6e78e2ca",
  1468 => x"d081c849",
  1469 => x"496e5166",
  1470 => x"66d481c9",
  1471 => x"ca496e51",
  1472 => x"5166dc81",
  1473 => x"c14866d0",
  1474 => x"58a6d480",
  1475 => x"cc4866c8",
  1476 => x"c004a866",
  1477 => x"66c887cb",
  1478 => x"cc80c148",
  1479 => x"d9c558a6",
  1480 => x"4866cc87",
  1481 => x"a6d088c1",
  1482 => x"87cec558",
  1483 => x"87f6d8ff",
  1484 => x"58a6e8c0",
  1485 => x"87eed8ff",
  1486 => x"58a6e0c0",
  1487 => x"05a8ecc0",
  1488 => x"dc87cac0",
  1489 => x"e4c048a6",
  1490 => x"c4c07866",
  1491 => x"e2d5ff87",
  1492 => x"4966c887",
  1493 => x"fcc091cb",
  1494 => x"80714866",
  1495 => x"c84a7e70",
  1496 => x"ca496e82",
  1497 => x"66e4c081",
  1498 => x"4966dc51",
  1499 => x"e4c081c1",
  1500 => x"48c18966",
  1501 => x"49703071",
  1502 => x"977189c1",
  1503 => x"c8f9c27a",
  1504 => x"e4c049bf",
  1505 => x"6a972966",
  1506 => x"9871484a",
  1507 => x"58a6ecc0",
  1508 => x"81c4496e",
  1509 => x"66d84d69",
  1510 => x"a866c448",
  1511 => x"87c8c002",
  1512 => x"c048a6c4",
  1513 => x"87c5c078",
  1514 => x"c148a6c4",
  1515 => x"1e66c478",
  1516 => x"751ee0c0",
  1517 => x"fed4ff49",
  1518 => x"7086c887",
  1519 => x"acb7c04c",
  1520 => x"87d4c106",
  1521 => x"e0c08574",
  1522 => x"75897449",
  1523 => x"f5e3c14b",
  1524 => x"e3fe714a",
  1525 => x"85c287d1",
  1526 => x"4866e0c0",
  1527 => x"e4c080c1",
  1528 => x"e8c058a6",
  1529 => x"81c14966",
  1530 => x"c002a970",
  1531 => x"a6c487c8",
  1532 => x"c078c048",
  1533 => x"a6c487c5",
  1534 => x"c478c148",
  1535 => x"a4c21e66",
  1536 => x"48e0c049",
  1537 => x"49708871",
  1538 => x"ff49751e",
  1539 => x"c887e8d3",
  1540 => x"a8b7c086",
  1541 => x"87c0ff01",
  1542 => x"0266e0c0",
  1543 => x"6e87d1c0",
  1544 => x"c081c949",
  1545 => x"6e5166e0",
  1546 => x"e3cbc148",
  1547 => x"87ccc078",
  1548 => x"81c9496e",
  1549 => x"486e51c2",
  1550 => x"78cfcdc1",
  1551 => x"cc4866c8",
  1552 => x"c004a866",
  1553 => x"66c887cb",
  1554 => x"cc80c148",
  1555 => x"e9c058a6",
  1556 => x"4866cc87",
  1557 => x"a6d088c1",
  1558 => x"87dec058",
  1559 => x"87c3d2ff",
  1560 => x"d5c04c70",
  1561 => x"acc6c187",
  1562 => x"87c8c005",
  1563 => x"c14866d0",
  1564 => x"58a6d480",
  1565 => x"87ebd1ff",
  1566 => x"66d44c70",
  1567 => x"d880c148",
  1568 => x"9c7458a6",
  1569 => x"87cbc002",
  1570 => x"c14866c8",
  1571 => x"04a866c4",
  1572 => x"ff87f7f2",
  1573 => x"c887c3d1",
  1574 => x"a8c74866",
  1575 => x"87e5c003",
  1576 => x"48dcf5c2",
  1577 => x"66c878c0",
  1578 => x"c091cb49",
  1579 => x"c48166fc",
  1580 => x"4a6a4aa1",
  1581 => x"c87952c0",
  1582 => x"80c14866",
  1583 => x"c758a6cc",
  1584 => x"dbff04a8",
  1585 => x"8ed4ff87",
  1586 => x"87e9dbff",
  1587 => x"64616f4c",
  1588 => x"74655320",
  1589 => x"676e6974",
  1590 => x"00812073",
  1591 => x"65766153",
  1592 => x"74655320",
  1593 => x"676e6974",
  1594 => x"00812073",
  1595 => x"64616f4c",
  1596 => x"202e2a20",
  1597 => x"00203a00",
  1598 => x"711e731e",
  1599 => x"c6029b4b",
  1600 => x"d8f5c287",
  1601 => x"c778c048",
  1602 => x"d8f5c21e",
  1603 => x"e8c11ebf",
  1604 => x"f5c21ec3",
  1605 => x"eb49bfc0",
  1606 => x"86cc87e4",
  1607 => x"bfc0f5c2",
  1608 => x"87cde049",
  1609 => x"c8029b73",
  1610 => x"c3e8c187",
  1611 => x"c8e2c049",
  1612 => x"c4daff87",
  1613 => x"c1c81e87",
  1614 => x"fe49c187",
  1615 => x"f5c287fa",
  1616 => x"50c048e0",
  1617 => x"87cfe6fe",
  1618 => x"cd029870",
  1619 => x"c9effe87",
  1620 => x"02987087",
  1621 => x"4ac187c4",
  1622 => x"4ac087c2",
  1623 => x"ce059a72",
  1624 => x"c11ec087",
  1625 => x"c049eae6",
  1626 => x"c487c5f2",
  1627 => x"c187fe86",
  1628 => x"c049f5e6",
  1629 => x"c287c7fc",
  1630 => x"c048d8f5",
  1631 => x"c0f5c278",
  1632 => x"1e78c048",
  1633 => x"49c1e7c1",
  1634 => x"87e4f1c0",
  1635 => x"ffc01ec0",
  1636 => x"497087d1",
  1637 => x"87d8f1c0",
  1638 => x"dcc386c8",
  1639 => x"dbe2c087",
  1640 => x"daf5c087",
  1641 => x"87f5ff87",
  1642 => x"44534f26",
  1643 => x"69616620",
  1644 => x"2e64656c",
  1645 => x"43495600",
  1646 => x"20203032",
  1647 => x"47464320",
  1648 => x"6f6f4200",
  1649 => x"676e6974",
  1650 => x"002e2e2e",
  1651 => x"00010000",
  1652 => x"20200000",
  1653 => x"20202020",
  1654 => x"20202020",
  1655 => x"45202020",
  1656 => x"20746978",
  1657 => x"20202020",
  1658 => x"20202020",
  1659 => x"81202020",
  1660 => x"20208000",
  1661 => x"20202020",
  1662 => x"20202020",
  1663 => x"61422020",
  1664 => x"5e006b63",
  1665 => x"6c000010",
  1666 => x"0000002d",
  1667 => x"105e0000",
  1668 => x"2d8a0000",
  1669 => x"00000000",
  1670 => x"00105e00",
  1671 => x"002da800",
  1672 => x"00000000",
  1673 => x"0000105e",
  1674 => x"00002dc6",
  1675 => x"5e000000",
  1676 => x"e4000010",
  1677 => x"0000002d",
  1678 => x"105e0000",
  1679 => x"2e020000",
  1680 => x"00000000",
  1681 => x"00105e00",
  1682 => x"002e2000",
  1683 => x"00000000",
  1684 => x"00001112",
  1685 => x"00000000",
  1686 => x"60000000",
  1687 => x"00000013",
  1688 => x"00000000",
  1689 => x"fe1e0000",
  1690 => x"78c048f0",
  1691 => x"097909cd",
  1692 => x"fe1e4f26",
  1693 => x"2648bff0",
  1694 => x"f0fe1e4f",
  1695 => x"2678c148",
  1696 => x"f0fe1e4f",
  1697 => x"2678c048",
  1698 => x"4a711e4f",
  1699 => x"265152c0",
  1700 => x"5b5e0e4f",
  1701 => x"f40e5d5c",
  1702 => x"974d7186",
  1703 => x"a5c17e6d",
  1704 => x"486c974c",
  1705 => x"6e58a6c8",
  1706 => x"a866c448",
  1707 => x"ff87c505",
  1708 => x"87e6c048",
  1709 => x"c287caff",
  1710 => x"6c9749a5",
  1711 => x"4ba3714b",
  1712 => x"974b6b97",
  1713 => x"486e7e6c",
  1714 => x"a6c880c1",
  1715 => x"cc98c758",
  1716 => x"977058a6",
  1717 => x"87e1fe7c",
  1718 => x"8ef44873",
  1719 => x"4c264d26",
  1720 => x"4f264b26",
  1721 => x"5c5b5e0e",
  1722 => x"7186f40e",
  1723 => x"4a66d84c",
  1724 => x"c29affc3",
  1725 => x"6c974ba4",
  1726 => x"49a17349",
  1727 => x"6c975172",
  1728 => x"c1486e7e",
  1729 => x"58a6c880",
  1730 => x"a6cc98c7",
  1731 => x"f4547058",
  1732 => x"87caff8e",
  1733 => x"e8fd1e1e",
  1734 => x"4abfe087",
  1735 => x"c0e0c049",
  1736 => x"87cb0299",
  1737 => x"f8c21e72",
  1738 => x"f7fe49fe",
  1739 => x"fd86c487",
  1740 => x"7e7087c0",
  1741 => x"2687c2fd",
  1742 => x"c21e4f26",
  1743 => x"fd49fef8",
  1744 => x"ecc187c7",
  1745 => x"ddfc49d4",
  1746 => x"87f5c287",
  1747 => x"731e4f26",
  1748 => x"fef8c21e",
  1749 => x"87f9fc49",
  1750 => x"b7c04a70",
  1751 => x"ccc204aa",
  1752 => x"aaf0c387",
  1753 => x"c187c905",
  1754 => x"c148f9ef",
  1755 => x"87edc178",
  1756 => x"05aae0c3",
  1757 => x"efc187c9",
  1758 => x"78c148fd",
  1759 => x"c187dec1",
  1760 => x"02bffdef",
  1761 => x"c0c287c6",
  1762 => x"87c24ba2",
  1763 => x"efc14b72",
  1764 => x"c002bff9",
  1765 => x"497387e0",
  1766 => x"9129b7c4",
  1767 => x"81d0f1c1",
  1768 => x"9acf4a73",
  1769 => x"48c192c2",
  1770 => x"4a703072",
  1771 => x"4872baff",
  1772 => x"79709869",
  1773 => x"497387db",
  1774 => x"9129b7c4",
  1775 => x"81d0f1c1",
  1776 => x"9acf4a73",
  1777 => x"48c392c2",
  1778 => x"4a703072",
  1779 => x"70b06948",
  1780 => x"fdefc179",
  1781 => x"c178c048",
  1782 => x"c048f9ef",
  1783 => x"fef8c278",
  1784 => x"87edfa49",
  1785 => x"b7c04a70",
  1786 => x"f4fd03aa",
  1787 => x"c448c087",
  1788 => x"264d2687",
  1789 => x"264b264c",
  1790 => x"0000004f",
  1791 => x"00000000",
  1792 => x"4ac01e00",
  1793 => x"91c44972",
  1794 => x"81d0f1c1",
  1795 => x"82c179c0",
  1796 => x"04aab7d0",
  1797 => x"4f2687ee",
  1798 => x"5c5b5e0e",
  1799 => x"4d710e5d",
  1800 => x"7587def9",
  1801 => x"2ab7c44a",
  1802 => x"d0f1c192",
  1803 => x"cf4c7582",
  1804 => x"6a94c29c",
  1805 => x"2b744b49",
  1806 => x"48c29bc3",
  1807 => x"4c703074",
  1808 => x"4874bcff",
  1809 => x"7a709871",
  1810 => x"7387eef8",
  1811 => x"87e1fe48",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"00000000",
  1817 => x"00000000",
  1818 => x"00000000",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"48d0ff1e",
  1829 => x"7178e1c8",
  1830 => x"08d4ff48",
  1831 => x"1e4f2678",
  1832 => x"c848d0ff",
  1833 => x"487178e1",
  1834 => x"7808d4ff",
  1835 => x"ff4866c4",
  1836 => x"267808d4",
  1837 => x"4a711e4f",
  1838 => x"1e4966c4",
  1839 => x"deff4972",
  1840 => x"48d0ff87",
  1841 => x"2678e0c0",
  1842 => x"731e4f26",
  1843 => x"c84b711e",
  1844 => x"731e4966",
  1845 => x"a2e0c14a",
  1846 => x"87d9ff49",
  1847 => x"2687c426",
  1848 => x"264c264d",
  1849 => x"1e4f264b",
  1850 => x"c34ad4ff",
  1851 => x"d0ff7aff",
  1852 => x"78e1c048",
  1853 => x"f9c27ade",
  1854 => x"497abfc8",
  1855 => x"7028c848",
  1856 => x"d048717a",
  1857 => x"717a7028",
  1858 => x"7028d848",
  1859 => x"48d0ff7a",
  1860 => x"2678e0c0",
  1861 => x"d0ff1e4f",
  1862 => x"78c9c848",
  1863 => x"d4ff4871",
  1864 => x"4f267808",
  1865 => x"494a711e",
  1866 => x"d0ff87eb",
  1867 => x"2678c848",
  1868 => x"1e731e4f",
  1869 => x"f9c24b71",
  1870 => x"c302bfd8",
  1871 => x"87ebc287",
  1872 => x"c848d0ff",
  1873 => x"487378c9",
  1874 => x"ffb0e0c0",
  1875 => x"c27808d4",
  1876 => x"c048ccf9",
  1877 => x"0266c878",
  1878 => x"ffc387c5",
  1879 => x"c087c249",
  1880 => x"d4f9c249",
  1881 => x"0266cc59",
  1882 => x"d5c587c6",
  1883 => x"87c44ad5",
  1884 => x"4affffcf",
  1885 => x"5ad8f9c2",
  1886 => x"48d8f9c2",
  1887 => x"87c478c1",
  1888 => x"4c264d26",
  1889 => x"4f264b26",
  1890 => x"5c5b5e0e",
  1891 => x"4a710e5d",
  1892 => x"bfd4f9c2",
  1893 => x"029a724c",
  1894 => x"c84987cb",
  1895 => x"e7f4c191",
  1896 => x"c483714b",
  1897 => x"e7f8c187",
  1898 => x"134dc04b",
  1899 => x"c2997449",
  1900 => x"48bfd0f9",
  1901 => x"d4ffb871",
  1902 => x"b7c17808",
  1903 => x"b7c8852c",
  1904 => x"87e704ad",
  1905 => x"bfccf9c2",
  1906 => x"c280c848",
  1907 => x"fe58d0f9",
  1908 => x"731e87ee",
  1909 => x"134b711e",
  1910 => x"cb029a4a",
  1911 => x"fe497287",
  1912 => x"4a1387e6",
  1913 => x"87f5059a",
  1914 => x"1e87d9fe",
  1915 => x"bfccf9c2",
  1916 => x"ccf9c249",
  1917 => x"78a1c148",
  1918 => x"a9b7c0c4",
  1919 => x"ff87db03",
  1920 => x"f9c248d4",
  1921 => x"c278bfd0",
  1922 => x"49bfccf9",
  1923 => x"48ccf9c2",
  1924 => x"c478a1c1",
  1925 => x"04a9b7c0",
  1926 => x"d0ff87e5",
  1927 => x"c278c848",
  1928 => x"c048d8f9",
  1929 => x"004f2678",
  1930 => x"00000000",
  1931 => x"00000000",
  1932 => x"5f5f0000",
  1933 => x"00000000",
  1934 => x"03000303",
  1935 => x"14000003",
  1936 => x"7f147f7f",
  1937 => x"0000147f",
  1938 => x"6b6b2e24",
  1939 => x"4c00123a",
  1940 => x"6c18366a",
  1941 => x"30003256",
  1942 => x"77594f7e",
  1943 => x"0040683a",
  1944 => x"03070400",
  1945 => x"00000000",
  1946 => x"633e1c00",
  1947 => x"00000041",
  1948 => x"3e634100",
  1949 => x"0800001c",
  1950 => x"1c1c3e2a",
  1951 => x"00082a3e",
  1952 => x"3e3e0808",
  1953 => x"00000808",
  1954 => x"60e08000",
  1955 => x"00000000",
  1956 => x"08080808",
  1957 => x"00000808",
  1958 => x"60600000",
  1959 => x"40000000",
  1960 => x"0c183060",
  1961 => x"00010306",
  1962 => x"4d597f3e",
  1963 => x"00003e7f",
  1964 => x"7f7f0604",
  1965 => x"00000000",
  1966 => x"59716342",
  1967 => x"0000464f",
  1968 => x"49496322",
  1969 => x"1800367f",
  1970 => x"7f13161c",
  1971 => x"0000107f",
  1972 => x"45456727",
  1973 => x"0000397d",
  1974 => x"494b7e3c",
  1975 => x"00003079",
  1976 => x"79710101",
  1977 => x"0000070f",
  1978 => x"49497f36",
  1979 => x"0000367f",
  1980 => x"69494f06",
  1981 => x"00001e3f",
  1982 => x"66660000",
  1983 => x"00000000",
  1984 => x"66e68000",
  1985 => x"00000000",
  1986 => x"14140808",
  1987 => x"00002222",
  1988 => x"14141414",
  1989 => x"00001414",
  1990 => x"14142222",
  1991 => x"00000808",
  1992 => x"59510302",
  1993 => x"3e00060f",
  1994 => x"555d417f",
  1995 => x"00001e1f",
  1996 => x"09097f7e",
  1997 => x"00007e7f",
  1998 => x"49497f7f",
  1999 => x"0000367f",
  2000 => x"41633e1c",
  2001 => x"00004141",
  2002 => x"63417f7f",
  2003 => x"00001c3e",
  2004 => x"49497f7f",
  2005 => x"00004141",
  2006 => x"09097f7f",
  2007 => x"00000101",
  2008 => x"49417f3e",
  2009 => x"00007a7b",
  2010 => x"08087f7f",
  2011 => x"00007f7f",
  2012 => x"7f7f4100",
  2013 => x"00000041",
  2014 => x"40406020",
  2015 => x"7f003f7f",
  2016 => x"361c087f",
  2017 => x"00004163",
  2018 => x"40407f7f",
  2019 => x"7f004040",
  2020 => x"060c067f",
  2021 => x"7f007f7f",
  2022 => x"180c067f",
  2023 => x"00007f7f",
  2024 => x"41417f3e",
  2025 => x"00003e7f",
  2026 => x"09097f7f",
  2027 => x"3e00060f",
  2028 => x"7f61417f",
  2029 => x"0000407e",
  2030 => x"19097f7f",
  2031 => x"0000667f",
  2032 => x"594d6f26",
  2033 => x"0000327b",
  2034 => x"7f7f0101",
  2035 => x"00000101",
  2036 => x"40407f3f",
  2037 => x"00003f7f",
  2038 => x"70703f0f",
  2039 => x"7f000f3f",
  2040 => x"3018307f",
  2041 => x"41007f7f",
  2042 => x"1c1c3663",
  2043 => x"01416336",
  2044 => x"7c7c0603",
  2045 => x"61010306",
  2046 => x"474d5971",
  2047 => x"00004143",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
