
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d4",x"ea",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"d4",x"ea",x"c2"),
    18 => (x"48",x"e4",x"d7",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"e4",x"d7",x"c2",x"87"),
    25 => (x"e0",x"d7",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e2",x"c1",x"87",x"f7"),
    29 => (x"d7",x"c2",x"87",x"d4"),
    30 => (x"d7",x"c2",x"4d",x"e4"),
    31 => (x"ad",x"74",x"4c",x"e4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"cf",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"df",x"4c",x"87",x"c9"),
    69 => (x"88",x"74",x"9c",x"98"),
    70 => (x"26",x"87",x"ec",x"02"),
    71 => (x"26",x"4b",x"26",x"4a"),
    72 => (x"1e",x"4f",x"26",x"4c"),
    73 => (x"73",x"81",x"48",x"73"),
    74 => (x"87",x"c5",x"02",x"a9"),
    75 => (x"f6",x"05",x"53",x"12"),
    76 => (x"0e",x"4f",x"26",x"87"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"d7",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"e4"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"e4",x"d7"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"e8",x"d7",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"c3",x"c3"),
   251 => (x"c2",x"58",x"ec",x"d7"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"fc",x"0e",x"5d",x"5c"),
   258 => (x"ff",x"4b",x"71",x"86"),
   259 => (x"7e",x"c0",x"4c",x"d4"),
   260 => (x"df",x"cd",x"ee",x"c5"),
   261 => (x"7c",x"ff",x"c3",x"4a"),
   262 => (x"fe",x"c3",x"48",x"6c"),
   263 => (x"f8",x"c0",x"05",x"a8"),
   264 => (x"73",x"4d",x"74",x"87"),
   265 => (x"87",x"cc",x"02",x"9b"),
   266 => (x"73",x"1e",x"66",x"d4"),
   267 => (x"87",x"c3",x"f4",x"49"),
   268 => (x"87",x"d4",x"86",x"c4"),
   269 => (x"c4",x"48",x"d0",x"ff"),
   270 => (x"66",x"d4",x"78",x"d1"),
   271 => (x"7d",x"ff",x"c3",x"4a"),
   272 => (x"f8",x"05",x"8a",x"c1"),
   273 => (x"5a",x"a6",x"d8",x"87"),
   274 => (x"7c",x"7c",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"4a",x"c1",x"78",x"d0"),
   278 => (x"05",x"8a",x"c1",x"7e"),
   279 => (x"6e",x"87",x"f6",x"fe"),
   280 => (x"26",x"8e",x"fc",x"48"),
   281 => (x"26",x"4c",x"26",x"4d"),
   282 => (x"1e",x"4f",x"26",x"4b"),
   283 => (x"4a",x"71",x"1e",x"73"),
   284 => (x"d4",x"ff",x"4b",x"c0"),
   285 => (x"78",x"ff",x"c3",x"48"),
   286 => (x"c4",x"48",x"d0",x"ff"),
   287 => (x"d4",x"ff",x"78",x"c3"),
   288 => (x"78",x"ff",x"c3",x"48"),
   289 => (x"ff",x"c0",x"1e",x"72"),
   290 => (x"49",x"d1",x"c1",x"f0"),
   291 => (x"c4",x"87",x"f9",x"f3"),
   292 => (x"05",x"98",x"70",x"86"),
   293 => (x"c0",x"c8",x"87",x"d2"),
   294 => (x"49",x"66",x"cc",x"1e"),
   295 => (x"c4",x"87",x"e2",x"fd"),
   296 => (x"ff",x"4b",x"70",x"86"),
   297 => (x"78",x"c2",x"48",x"d0"),
   298 => (x"4b",x"26",x"48",x"73"),
   299 => (x"5e",x"0e",x"4f",x"26"),
   300 => (x"0e",x"5d",x"5c",x"5b"),
   301 => (x"ff",x"c0",x"1e",x"c0"),
   302 => (x"49",x"c9",x"c1",x"f0"),
   303 => (x"d2",x"87",x"c9",x"f3"),
   304 => (x"f4",x"d7",x"c2",x"1e"),
   305 => (x"87",x"f9",x"fc",x"49"),
   306 => (x"4c",x"c0",x"86",x"c8"),
   307 => (x"b7",x"d2",x"84",x"c1"),
   308 => (x"87",x"f8",x"04",x"ac"),
   309 => (x"97",x"f4",x"d7",x"c2"),
   310 => (x"c0",x"c3",x"49",x"bf"),
   311 => (x"a9",x"c0",x"c1",x"99"),
   312 => (x"87",x"e7",x"c0",x"05"),
   313 => (x"97",x"fb",x"d7",x"c2"),
   314 => (x"31",x"d0",x"49",x"bf"),
   315 => (x"97",x"fc",x"d7",x"c2"),
   316 => (x"32",x"c8",x"4a",x"bf"),
   317 => (x"d7",x"c2",x"b1",x"72"),
   318 => (x"4a",x"bf",x"97",x"fd"),
   319 => (x"cf",x"4c",x"71",x"b1"),
   320 => (x"9c",x"ff",x"ff",x"ff"),
   321 => (x"34",x"ca",x"84",x"c1"),
   322 => (x"c2",x"87",x"e7",x"c1"),
   323 => (x"bf",x"97",x"fd",x"d7"),
   324 => (x"c6",x"31",x"c1",x"49"),
   325 => (x"fe",x"d7",x"c2",x"99"),
   326 => (x"c7",x"4a",x"bf",x"97"),
   327 => (x"b1",x"72",x"2a",x"b7"),
   328 => (x"97",x"f9",x"d7",x"c2"),
   329 => (x"cf",x"4d",x"4a",x"bf"),
   330 => (x"fa",x"d7",x"c2",x"9d"),
   331 => (x"c3",x"4a",x"bf",x"97"),
   332 => (x"c2",x"32",x"ca",x"9a"),
   333 => (x"bf",x"97",x"fb",x"d7"),
   334 => (x"73",x"33",x"c2",x"4b"),
   335 => (x"fc",x"d7",x"c2",x"b2"),
   336 => (x"c3",x"4b",x"bf",x"97"),
   337 => (x"b7",x"c6",x"9b",x"c0"),
   338 => (x"c2",x"b2",x"73",x"2b"),
   339 => (x"71",x"48",x"c1",x"81"),
   340 => (x"c1",x"49",x"70",x"30"),
   341 => (x"70",x"30",x"75",x"48"),
   342 => (x"c1",x"4c",x"72",x"4d"),
   343 => (x"c8",x"94",x"71",x"84"),
   344 => (x"06",x"ad",x"b7",x"c0"),
   345 => (x"34",x"c1",x"87",x"cc"),
   346 => (x"c0",x"c8",x"2d",x"b7"),
   347 => (x"ff",x"01",x"ad",x"b7"),
   348 => (x"48",x"74",x"87",x"f4"),
   349 => (x"4c",x"26",x"4d",x"26"),
   350 => (x"4f",x"26",x"4b",x"26"),
   351 => (x"5c",x"5b",x"5e",x"0e"),
   352 => (x"86",x"f8",x"0e",x"5d"),
   353 => (x"48",x"dc",x"e0",x"c2"),
   354 => (x"d8",x"c2",x"78",x"c0"),
   355 => (x"49",x"c0",x"1e",x"d4"),
   356 => (x"c4",x"87",x"d8",x"fb"),
   357 => (x"05",x"98",x"70",x"86"),
   358 => (x"48",x"c0",x"87",x"c5"),
   359 => (x"c0",x"87",x"f1",x"c8"),
   360 => (x"c2",x"7e",x"c1",x"4d"),
   361 => (x"df",x"4a",x"ca",x"d9"),
   362 => (x"4b",x"c8",x"49",x"e8"),
   363 => (x"70",x"87",x"f7",x"ec"),
   364 => (x"87",x"c2",x"05",x"98"),
   365 => (x"d9",x"c2",x"7e",x"c0"),
   366 => (x"f4",x"df",x"4a",x"e6"),
   367 => (x"ec",x"4b",x"c8",x"49"),
   368 => (x"98",x"70",x"87",x"e4"),
   369 => (x"c0",x"87",x"c2",x"05"),
   370 => (x"c0",x"02",x"6e",x"7e"),
   371 => (x"df",x"c2",x"87",x"fd"),
   372 => (x"c2",x"4d",x"bf",x"da"),
   373 => (x"bf",x"9f",x"d2",x"e0"),
   374 => (x"d6",x"c5",x"48",x"7e"),
   375 => (x"c7",x"05",x"a8",x"ea"),
   376 => (x"da",x"df",x"c2",x"87"),
   377 => (x"87",x"ce",x"4d",x"bf"),
   378 => (x"e9",x"ca",x"48",x"6e"),
   379 => (x"c5",x"02",x"a8",x"d5"),
   380 => (x"c7",x"48",x"c0",x"87"),
   381 => (x"d8",x"c2",x"87",x"da"),
   382 => (x"49",x"75",x"1e",x"d4"),
   383 => (x"c4",x"87",x"ec",x"f9"),
   384 => (x"05",x"98",x"70",x"86"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c5",x"c7"),
   387 => (x"c0",x"4a",x"e6",x"d9"),
   388 => (x"c8",x"49",x"c0",x"e0"),
   389 => (x"87",x"ce",x"eb",x"4b"),
   390 => (x"c8",x"05",x"98",x"70"),
   391 => (x"dc",x"e0",x"c2",x"87"),
   392 => (x"d7",x"78",x"c1",x"48"),
   393 => (x"ca",x"d9",x"c2",x"87"),
   394 => (x"cc",x"e0",x"c0",x"4a"),
   395 => (x"ea",x"4b",x"c8",x"49"),
   396 => (x"98",x"70",x"87",x"f4"),
   397 => (x"c0",x"87",x"c5",x"02"),
   398 => (x"87",x"d4",x"c6",x"48"),
   399 => (x"97",x"d2",x"e0",x"c2"),
   400 => (x"d5",x"c1",x"49",x"bf"),
   401 => (x"87",x"cd",x"05",x"a9"),
   402 => (x"97",x"d3",x"e0",x"c2"),
   403 => (x"ea",x"c2",x"49",x"bf"),
   404 => (x"c5",x"c0",x"02",x"a9"),
   405 => (x"c5",x"48",x"c0",x"87"),
   406 => (x"d8",x"c2",x"87",x"f6"),
   407 => (x"7e",x"bf",x"97",x"d4"),
   408 => (x"a8",x"e9",x"c3",x"48"),
   409 => (x"87",x"ce",x"c0",x"02"),
   410 => (x"eb",x"c3",x"48",x"6e"),
   411 => (x"c5",x"c0",x"02",x"a8"),
   412 => (x"c5",x"48",x"c0",x"87"),
   413 => (x"d8",x"c2",x"87",x"da"),
   414 => (x"49",x"bf",x"97",x"df"),
   415 => (x"cc",x"c0",x"05",x"99"),
   416 => (x"e0",x"d8",x"c2",x"87"),
   417 => (x"c2",x"49",x"bf",x"97"),
   418 => (x"c5",x"c0",x"02",x"a9"),
   419 => (x"c4",x"48",x"c0",x"87"),
   420 => (x"d8",x"c2",x"87",x"fe"),
   421 => (x"48",x"bf",x"97",x"e1"),
   422 => (x"58",x"d8",x"e0",x"c2"),
   423 => (x"c1",x"48",x"4c",x"70"),
   424 => (x"dc",x"e0",x"c2",x"88"),
   425 => (x"e2",x"d8",x"c2",x"58"),
   426 => (x"75",x"49",x"bf",x"97"),
   427 => (x"e3",x"d8",x"c2",x"81"),
   428 => (x"c8",x"4a",x"bf",x"97"),
   429 => (x"7e",x"a1",x"72",x"32"),
   430 => (x"48",x"ec",x"e4",x"c2"),
   431 => (x"d8",x"c2",x"78",x"6e"),
   432 => (x"48",x"bf",x"97",x"e4"),
   433 => (x"c2",x"58",x"a6",x"c8"),
   434 => (x"02",x"bf",x"dc",x"e0"),
   435 => (x"c2",x"87",x"cc",x"c2"),
   436 => (x"df",x"4a",x"e6",x"d9"),
   437 => (x"4b",x"c8",x"49",x"dc"),
   438 => (x"70",x"87",x"cb",x"e8"),
   439 => (x"c5",x"c0",x"02",x"98"),
   440 => (x"c3",x"48",x"c0",x"87"),
   441 => (x"e0",x"c2",x"87",x"ea"),
   442 => (x"c2",x"4c",x"bf",x"d4"),
   443 => (x"c2",x"5c",x"c0",x"e5"),
   444 => (x"bf",x"97",x"f9",x"d8"),
   445 => (x"c2",x"31",x"c8",x"49"),
   446 => (x"bf",x"97",x"f8",x"d8"),
   447 => (x"c2",x"49",x"a1",x"4a"),
   448 => (x"bf",x"97",x"fa",x"d8"),
   449 => (x"72",x"32",x"d0",x"4a"),
   450 => (x"d8",x"c2",x"49",x"a1"),
   451 => (x"4a",x"bf",x"97",x"fb"),
   452 => (x"a1",x"72",x"32",x"d8"),
   453 => (x"91",x"66",x"c4",x"49"),
   454 => (x"bf",x"ec",x"e4",x"c2"),
   455 => (x"f4",x"e4",x"c2",x"81"),
   456 => (x"c1",x"d9",x"c2",x"59"),
   457 => (x"c8",x"4a",x"bf",x"97"),
   458 => (x"c0",x"d9",x"c2",x"32"),
   459 => (x"a2",x"4b",x"bf",x"97"),
   460 => (x"c2",x"d9",x"c2",x"4a"),
   461 => (x"d0",x"4b",x"bf",x"97"),
   462 => (x"4a",x"a2",x"73",x"33"),
   463 => (x"97",x"c3",x"d9",x"c2"),
   464 => (x"9b",x"cf",x"4b",x"bf"),
   465 => (x"a2",x"73",x"33",x"d8"),
   466 => (x"f8",x"e4",x"c2",x"4a"),
   467 => (x"74",x"8a",x"c2",x"5a"),
   468 => (x"f8",x"e4",x"c2",x"92"),
   469 => (x"78",x"a1",x"72",x"48"),
   470 => (x"c2",x"87",x"c1",x"c1"),
   471 => (x"bf",x"97",x"e6",x"d8"),
   472 => (x"c2",x"31",x"c8",x"49"),
   473 => (x"bf",x"97",x"e5",x"d8"),
   474 => (x"c5",x"49",x"a1",x"4a"),
   475 => (x"81",x"ff",x"c7",x"31"),
   476 => (x"e5",x"c2",x"29",x"c9"),
   477 => (x"d8",x"c2",x"59",x"c0"),
   478 => (x"4a",x"bf",x"97",x"eb"),
   479 => (x"d8",x"c2",x"32",x"c8"),
   480 => (x"4b",x"bf",x"97",x"ea"),
   481 => (x"66",x"c4",x"4a",x"a2"),
   482 => (x"c2",x"82",x"6e",x"92"),
   483 => (x"c2",x"5a",x"fc",x"e4"),
   484 => (x"c0",x"48",x"f4",x"e4"),
   485 => (x"f0",x"e4",x"c2",x"78"),
   486 => (x"78",x"a1",x"72",x"48"),
   487 => (x"48",x"c0",x"e5",x"c2"),
   488 => (x"bf",x"f4",x"e4",x"c2"),
   489 => (x"c4",x"e5",x"c2",x"78"),
   490 => (x"f8",x"e4",x"c2",x"48"),
   491 => (x"e0",x"c2",x"78",x"bf"),
   492 => (x"c0",x"02",x"bf",x"dc"),
   493 => (x"48",x"74",x"87",x"c9"),
   494 => (x"7e",x"70",x"30",x"c4"),
   495 => (x"c2",x"87",x"c9",x"c0"),
   496 => (x"48",x"bf",x"fc",x"e4"),
   497 => (x"7e",x"70",x"30",x"c4"),
   498 => (x"48",x"e0",x"e0",x"c2"),
   499 => (x"48",x"c1",x"78",x"6e"),
   500 => (x"4d",x"26",x"8e",x"f8"),
   501 => (x"4b",x"26",x"4c",x"26"),
   502 => (x"00",x"00",x"4f",x"26"),
   503 => (x"33",x"54",x"41",x"46"),
   504 => (x"20",x"20",x"20",x"32"),
   505 => (x"00",x"00",x"00",x"00"),
   506 => (x"31",x"54",x"41",x"46"),
   507 => (x"20",x"20",x"20",x"36"),
   508 => (x"00",x"00",x"00",x"00"),
   509 => (x"33",x"54",x"41",x"46"),
   510 => (x"20",x"20",x"20",x"32"),
   511 => (x"00",x"00",x"00",x"00"),
   512 => (x"33",x"54",x"41",x"46"),
   513 => (x"20",x"20",x"20",x"32"),
   514 => (x"00",x"00",x"00",x"00"),
   515 => (x"31",x"54",x"41",x"46"),
   516 => (x"20",x"20",x"20",x"36"),
   517 => (x"00",x"00",x"00",x"00"),
   518 => (x"20",x"20",x"2e",x"2e"),
   519 => (x"20",x"20",x"20",x"20"),
   520 => (x"00",x"20",x"20",x"20"),
   521 => (x"5c",x"5b",x"5e",x"0e"),
   522 => (x"4a",x"71",x"0e",x"5d"),
   523 => (x"bf",x"dc",x"e0",x"c2"),
   524 => (x"72",x"87",x"cb",x"02"),
   525 => (x"72",x"2b",x"c7",x"4b"),
   526 => (x"9d",x"ff",x"c1",x"4d"),
   527 => (x"4b",x"72",x"87",x"c9"),
   528 => (x"4d",x"72",x"2b",x"c8"),
   529 => (x"c2",x"9d",x"ff",x"c3"),
   530 => (x"83",x"bf",x"ec",x"e4"),
   531 => (x"bf",x"d4",x"f2",x"c0"),
   532 => (x"87",x"d9",x"02",x"ab"),
   533 => (x"5b",x"d8",x"f2",x"c0"),
   534 => (x"1e",x"d4",x"d8",x"c2"),
   535 => (x"ca",x"f0",x"49",x"73"),
   536 => (x"70",x"86",x"c4",x"87"),
   537 => (x"87",x"c5",x"05",x"98"),
   538 => (x"e6",x"c0",x"48",x"c0"),
   539 => (x"dc",x"e0",x"c2",x"87"),
   540 => (x"87",x"d2",x"02",x"bf"),
   541 => (x"91",x"c4",x"49",x"75"),
   542 => (x"81",x"d4",x"d8",x"c2"),
   543 => (x"ff",x"cf",x"4c",x"69"),
   544 => (x"9c",x"ff",x"ff",x"ff"),
   545 => (x"49",x"75",x"87",x"cb"),
   546 => (x"d8",x"c2",x"91",x"c2"),
   547 => (x"69",x"9f",x"81",x"d4"),
   548 => (x"26",x"48",x"74",x"4c"),
   549 => (x"26",x"4c",x"26",x"4d"),
   550 => (x"0e",x"4f",x"26",x"4b"),
   551 => (x"5d",x"5c",x"5b",x"5e"),
   552 => (x"cc",x"86",x"f4",x"0e"),
   553 => (x"66",x"dc",x"59",x"a6"),
   554 => (x"dc",x"87",x"c7",x"02"),
   555 => (x"05",x"bf",x"97",x"66"),
   556 => (x"48",x"c0",x"87",x"c5"),
   557 => (x"c8",x"87",x"f4",x"c2"),
   558 => (x"80",x"c8",x"48",x"66"),
   559 => (x"c0",x"48",x"7e",x"70"),
   560 => (x"49",x"c1",x"1e",x"78"),
   561 => (x"87",x"d4",x"c7",x"49"),
   562 => (x"4c",x"70",x"86",x"c4"),
   563 => (x"fb",x"c0",x"02",x"9c"),
   564 => (x"e4",x"e0",x"c2",x"87"),
   565 => (x"49",x"66",x"dc",x"4a"),
   566 => (x"87",x"ef",x"df",x"ff"),
   567 => (x"c0",x"02",x"98",x"70"),
   568 => (x"4a",x"74",x"87",x"ea"),
   569 => (x"cb",x"49",x"66",x"dc"),
   570 => (x"87",x"d4",x"e0",x"4b"),
   571 => (x"db",x"02",x"98",x"70"),
   572 => (x"74",x"1e",x"c0",x"87"),
   573 => (x"87",x"c4",x"02",x"9c"),
   574 => (x"87",x"c2",x"4d",x"c0"),
   575 => (x"49",x"75",x"4d",x"c1"),
   576 => (x"c4",x"87",x"d9",x"c6"),
   577 => (x"9c",x"4c",x"70",x"86"),
   578 => (x"87",x"c5",x"ff",x"05"),
   579 => (x"c1",x"02",x"9c",x"74"),
   580 => (x"a4",x"dc",x"87",x"d7"),
   581 => (x"69",x"48",x"6e",x"49"),
   582 => (x"49",x"a4",x"da",x"78"),
   583 => (x"c4",x"48",x"66",x"c8"),
   584 => (x"58",x"a6",x"c8",x"80"),
   585 => (x"c4",x"48",x"69",x"9f"),
   586 => (x"c2",x"78",x"08",x"66"),
   587 => (x"02",x"bf",x"dc",x"e0"),
   588 => (x"a4",x"d4",x"87",x"d2"),
   589 => (x"49",x"69",x"9f",x"49"),
   590 => (x"99",x"ff",x"ff",x"c0"),
   591 => (x"30",x"d0",x"48",x"71"),
   592 => (x"87",x"c2",x"7e",x"70"),
   593 => (x"48",x"6e",x"7e",x"c0"),
   594 => (x"80",x"bf",x"66",x"c4"),
   595 => (x"78",x"08",x"66",x"c4"),
   596 => (x"c0",x"48",x"66",x"c8"),
   597 => (x"49",x"66",x"c8",x"78"),
   598 => (x"66",x"c4",x"81",x"cc"),
   599 => (x"66",x"c8",x"79",x"bf"),
   600 => (x"c0",x"81",x"d0",x"49"),
   601 => (x"c2",x"48",x"c1",x"79"),
   602 => (x"f4",x"48",x"c0",x"87"),
   603 => (x"26",x"4d",x"26",x"8e"),
   604 => (x"26",x"4b",x"26",x"4c"),
   605 => (x"5b",x"5e",x"0e",x"4f"),
   606 => (x"71",x"0e",x"5d",x"5c"),
   607 => (x"4d",x"66",x"d0",x"4c"),
   608 => (x"72",x"49",x"6c",x"4a"),
   609 => (x"c2",x"b9",x"4d",x"a1"),
   610 => (x"4a",x"bf",x"d8",x"e0"),
   611 => (x"99",x"72",x"ba",x"ff"),
   612 => (x"c0",x"02",x"99",x"71"),
   613 => (x"a4",x"c4",x"87",x"e4"),
   614 => (x"fa",x"49",x"6b",x"4b"),
   615 => (x"7b",x"70",x"87",x"c6"),
   616 => (x"bf",x"d4",x"e0",x"c2"),
   617 => (x"71",x"81",x"6c",x"49"),
   618 => (x"c2",x"b9",x"75",x"7c"),
   619 => (x"4a",x"bf",x"d8",x"e0"),
   620 => (x"99",x"72",x"ba",x"ff"),
   621 => (x"ff",x"05",x"99",x"71"),
   622 => (x"7c",x"75",x"87",x"dc"),
   623 => (x"4c",x"26",x"4d",x"26"),
   624 => (x"4f",x"26",x"4b",x"26"),
   625 => (x"71",x"1e",x"73",x"1e"),
   626 => (x"f0",x"e4",x"c2",x"4b"),
   627 => (x"a3",x"c4",x"49",x"bf"),
   628 => (x"c2",x"4a",x"6a",x"4a"),
   629 => (x"d4",x"e0",x"c2",x"8a"),
   630 => (x"a1",x"72",x"92",x"bf"),
   631 => (x"d8",x"e0",x"c2",x"49"),
   632 => (x"9a",x"6b",x"4a",x"bf"),
   633 => (x"c0",x"49",x"a1",x"72"),
   634 => (x"c8",x"59",x"d8",x"f2"),
   635 => (x"e9",x"71",x"1e",x"66"),
   636 => (x"86",x"c4",x"87",x"f9"),
   637 => (x"c4",x"05",x"98",x"70"),
   638 => (x"c2",x"48",x"c0",x"87"),
   639 => (x"26",x"48",x"c1",x"87"),
   640 => (x"1e",x"4f",x"26",x"4b"),
   641 => (x"4b",x"71",x"1e",x"73"),
   642 => (x"e4",x"c0",x"02",x"9b"),
   643 => (x"c4",x"e5",x"c2",x"87"),
   644 => (x"c2",x"4a",x"73",x"5b"),
   645 => (x"d4",x"e0",x"c2",x"8a"),
   646 => (x"c2",x"92",x"49",x"bf"),
   647 => (x"48",x"bf",x"f0",x"e4"),
   648 => (x"e5",x"c2",x"80",x"72"),
   649 => (x"48",x"71",x"58",x"c8"),
   650 => (x"e0",x"c2",x"30",x"c4"),
   651 => (x"ed",x"c0",x"58",x"e4"),
   652 => (x"c0",x"e5",x"c2",x"87"),
   653 => (x"f4",x"e4",x"c2",x"48"),
   654 => (x"e5",x"c2",x"78",x"bf"),
   655 => (x"e4",x"c2",x"48",x"c4"),
   656 => (x"c2",x"78",x"bf",x"f8"),
   657 => (x"02",x"bf",x"dc",x"e0"),
   658 => (x"e0",x"c2",x"87",x"c9"),
   659 => (x"c4",x"49",x"bf",x"d4"),
   660 => (x"c2",x"87",x"c7",x"31"),
   661 => (x"49",x"bf",x"fc",x"e4"),
   662 => (x"e0",x"c2",x"31",x"c4"),
   663 => (x"4b",x"26",x"59",x"e4"),
   664 => (x"5e",x"0e",x"4f",x"26"),
   665 => (x"71",x"0e",x"5c",x"5b"),
   666 => (x"72",x"4b",x"c0",x"4a"),
   667 => (x"e0",x"c0",x"02",x"9a"),
   668 => (x"49",x"a2",x"da",x"87"),
   669 => (x"c2",x"4b",x"69",x"9f"),
   670 => (x"02",x"bf",x"dc",x"e0"),
   671 => (x"a2",x"d4",x"87",x"cf"),
   672 => (x"49",x"69",x"9f",x"49"),
   673 => (x"ff",x"ff",x"c0",x"4c"),
   674 => (x"c2",x"34",x"d0",x"9c"),
   675 => (x"74",x"4c",x"c0",x"87"),
   676 => (x"fd",x"49",x"73",x"b3"),
   677 => (x"4c",x"26",x"87",x"ed"),
   678 => (x"4f",x"26",x"4b",x"26"),
   679 => (x"5c",x"5b",x"5e",x"0e"),
   680 => (x"86",x"f0",x"0e",x"5d"),
   681 => (x"cf",x"59",x"a6",x"c8"),
   682 => (x"f8",x"ff",x"ff",x"ff"),
   683 => (x"c4",x"7e",x"c0",x"4c"),
   684 => (x"87",x"d8",x"02",x"66"),
   685 => (x"48",x"d0",x"d8",x"c2"),
   686 => (x"d8",x"c2",x"78",x"c0"),
   687 => (x"e5",x"c2",x"48",x"c8"),
   688 => (x"c2",x"78",x"bf",x"c4"),
   689 => (x"c2",x"48",x"cc",x"d8"),
   690 => (x"78",x"bf",x"c0",x"e5"),
   691 => (x"48",x"f1",x"e0",x"c2"),
   692 => (x"e0",x"c2",x"50",x"c0"),
   693 => (x"c2",x"49",x"bf",x"e0"),
   694 => (x"4a",x"bf",x"d0",x"d8"),
   695 => (x"c4",x"03",x"aa",x"71"),
   696 => (x"49",x"72",x"87",x"cb"),
   697 => (x"c0",x"05",x"99",x"cf"),
   698 => (x"f2",x"c0",x"87",x"e9"),
   699 => (x"d8",x"c2",x"48",x"d4"),
   700 => (x"c2",x"78",x"bf",x"c8"),
   701 => (x"c2",x"1e",x"d4",x"d8"),
   702 => (x"49",x"bf",x"c8",x"d8"),
   703 => (x"48",x"c8",x"d8",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"e4",x"e5"),
   706 => (x"d0",x"f2",x"c0",x"86"),
   707 => (x"d4",x"d8",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"d0",x"f2"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"d4",x"f2"),
   712 => (x"48",x"bf",x"d0",x"d8"),
   713 => (x"d8",x"c2",x"80",x"c1"),
   714 => (x"90",x"27",x"58",x"d4"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e5",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"de",x"c2"),
   720 => (x"4b",x"bf",x"d0",x"f2"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"e4",x"e0"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"fc",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ed",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d3",x"05",x"99"),
   748 => (x"02",x"66",x"e0",x"c0"),
   749 => (x"73",x"87",x"cc",x"c0"),
   750 => (x"66",x"e0",x"c0",x"49"),
   751 => (x"02",x"98",x"70",x"0f"),
   752 => (x"6e",x"87",x"d3",x"c0"),
   753 => (x"87",x"c6",x"c0",x"05"),
   754 => (x"48",x"e4",x"e0",x"c2"),
   755 => (x"f2",x"c0",x"50",x"c0"),
   756 => (x"c2",x"48",x"bf",x"d0"),
   757 => (x"e0",x"c2",x"87",x"e9"),
   758 => (x"50",x"c0",x"48",x"f1"),
   759 => (x"e0",x"e0",x"c2",x"7e"),
   760 => (x"d8",x"c2",x"49",x"bf"),
   761 => (x"71",x"4a",x"bf",x"d0"),
   762 => (x"f5",x"fb",x"04",x"aa"),
   763 => (x"ff",x"ff",x"cf",x"87"),
   764 => (x"c2",x"4c",x"f8",x"ff"),
   765 => (x"05",x"bf",x"c4",x"e5"),
   766 => (x"c2",x"87",x"c8",x"c0"),
   767 => (x"02",x"bf",x"dc",x"e0"),
   768 => (x"c2",x"87",x"fa",x"c1"),
   769 => (x"49",x"bf",x"cc",x"d8"),
   770 => (x"c2",x"87",x"d9",x"f0"),
   771 => (x"c4",x"58",x"d0",x"d8"),
   772 => (x"d8",x"c2",x"48",x"a6"),
   773 => (x"c2",x"78",x"bf",x"cc"),
   774 => (x"02",x"bf",x"dc",x"e0"),
   775 => (x"c4",x"87",x"db",x"c0"),
   776 => (x"99",x"74",x"49",x"66"),
   777 => (x"c0",x"02",x"a9",x"74"),
   778 => (x"a6",x"c8",x"87",x"c8"),
   779 => (x"c0",x"78",x"c0",x"48"),
   780 => (x"a6",x"c8",x"87",x"e7"),
   781 => (x"c0",x"78",x"c1",x"48"),
   782 => (x"66",x"c4",x"87",x"df"),
   783 => (x"f8",x"ff",x"cf",x"49"),
   784 => (x"c0",x"02",x"a9",x"99"),
   785 => (x"a6",x"cc",x"87",x"c8"),
   786 => (x"c0",x"78",x"c0",x"48"),
   787 => (x"a6",x"cc",x"87",x"c5"),
   788 => (x"c8",x"78",x"c1",x"48"),
   789 => (x"66",x"cc",x"48",x"a6"),
   790 => (x"05",x"66",x"c8",x"78"),
   791 => (x"c4",x"87",x"de",x"c0"),
   792 => (x"89",x"c2",x"49",x"66"),
   793 => (x"bf",x"d4",x"e0",x"c2"),
   794 => (x"f0",x"e4",x"c2",x"91"),
   795 => (x"80",x"71",x"48",x"bf"),
   796 => (x"58",x"cc",x"d8",x"c2"),
   797 => (x"48",x"d0",x"d8",x"c2"),
   798 => (x"d5",x"f9",x"78",x"c0"),
   799 => (x"cf",x"48",x"c0",x"87"),
   800 => (x"f8",x"ff",x"ff",x"ff"),
   801 => (x"26",x"8e",x"f0",x"4c"),
   802 => (x"26",x"4c",x"26",x"4d"),
   803 => (x"00",x"4f",x"26",x"4b"),
   804 => (x"00",x"00",x"00",x"00"),
   805 => (x"ff",x"ff",x"ff",x"ff"),
   806 => (x"48",x"d4",x"ff",x"1e"),
   807 => (x"68",x"78",x"ff",x"c3"),
   808 => (x"1e",x"4f",x"26",x"48"),
   809 => (x"c3",x"48",x"d4",x"ff"),
   810 => (x"d0",x"ff",x"78",x"ff"),
   811 => (x"78",x"e1",x"c0",x"48"),
   812 => (x"d4",x"48",x"d4",x"ff"),
   813 => (x"1e",x"4f",x"26",x"78"),
   814 => (x"c0",x"48",x"d0",x"ff"),
   815 => (x"4f",x"26",x"78",x"e0"),
   816 => (x"87",x"d4",x"ff",x"1e"),
   817 => (x"02",x"99",x"49",x"70"),
   818 => (x"fb",x"c0",x"87",x"c6"),
   819 => (x"87",x"f1",x"05",x"a9"),
   820 => (x"4f",x"26",x"48",x"71"),
   821 => (x"5c",x"5b",x"5e",x"0e"),
   822 => (x"c0",x"4b",x"71",x"0e"),
   823 => (x"87",x"f8",x"fe",x"4c"),
   824 => (x"02",x"99",x"49",x"70"),
   825 => (x"c0",x"87",x"f9",x"c0"),
   826 => (x"c0",x"02",x"a9",x"ec"),
   827 => (x"fb",x"c0",x"87",x"f2"),
   828 => (x"eb",x"c0",x"02",x"a9"),
   829 => (x"b7",x"66",x"cc",x"87"),
   830 => (x"87",x"c7",x"03",x"ac"),
   831 => (x"c2",x"02",x"66",x"d0"),
   832 => (x"71",x"53",x"71",x"87"),
   833 => (x"87",x"c2",x"02",x"99"),
   834 => (x"cb",x"fe",x"84",x"c1"),
   835 => (x"99",x"49",x"70",x"87"),
   836 => (x"c0",x"87",x"cd",x"02"),
   837 => (x"c7",x"02",x"a9",x"ec"),
   838 => (x"a9",x"fb",x"c0",x"87"),
   839 => (x"87",x"d5",x"ff",x"05"),
   840 => (x"c3",x"02",x"66",x"d0"),
   841 => (x"7b",x"97",x"c0",x"87"),
   842 => (x"05",x"a9",x"ec",x"c0"),
   843 => (x"4a",x"74",x"87",x"c4"),
   844 => (x"4a",x"74",x"87",x"c5"),
   845 => (x"72",x"8a",x"0a",x"c0"),
   846 => (x"26",x"4c",x"26",x"48"),
   847 => (x"1e",x"4f",x"26",x"4b"),
   848 => (x"70",x"87",x"d5",x"fd"),
   849 => (x"f0",x"c0",x"4a",x"49"),
   850 => (x"87",x"c9",x"04",x"aa"),
   851 => (x"01",x"aa",x"f9",x"c0"),
   852 => (x"f0",x"c0",x"87",x"c3"),
   853 => (x"aa",x"c1",x"c1",x"8a"),
   854 => (x"c1",x"87",x"c9",x"04"),
   855 => (x"c3",x"01",x"aa",x"da"),
   856 => (x"8a",x"f7",x"c0",x"87"),
   857 => (x"4f",x"26",x"48",x"72"),
   858 => (x"5c",x"5b",x"5e",x"0e"),
   859 => (x"86",x"f8",x"0e",x"5d"),
   860 => (x"7e",x"c0",x"4c",x"71"),
   861 => (x"c0",x"87",x"ec",x"fc"),
   862 => (x"c8",x"f8",x"c0",x"4b"),
   863 => (x"c0",x"49",x"bf",x"97"),
   864 => (x"87",x"cf",x"04",x"a9"),
   865 => (x"c1",x"87",x"f9",x"fc"),
   866 => (x"c8",x"f8",x"c0",x"83"),
   867 => (x"ab",x"49",x"bf",x"97"),
   868 => (x"c0",x"87",x"f1",x"06"),
   869 => (x"bf",x"97",x"c8",x"f8"),
   870 => (x"fb",x"87",x"cf",x"02"),
   871 => (x"49",x"70",x"87",x"fa"),
   872 => (x"87",x"c6",x"02",x"99"),
   873 => (x"05",x"a9",x"ec",x"c0"),
   874 => (x"4b",x"c0",x"87",x"f1"),
   875 => (x"70",x"87",x"e9",x"fb"),
   876 => (x"87",x"e4",x"fb",x"4d"),
   877 => (x"fb",x"58",x"a6",x"c8"),
   878 => (x"4a",x"70",x"87",x"de"),
   879 => (x"a4",x"c8",x"83",x"c1"),
   880 => (x"49",x"69",x"97",x"49"),
   881 => (x"87",x"da",x"05",x"ad"),
   882 => (x"97",x"49",x"a4",x"c9"),
   883 => (x"66",x"c4",x"49",x"69"),
   884 => (x"87",x"ce",x"05",x"a9"),
   885 => (x"97",x"49",x"a4",x"ca"),
   886 => (x"05",x"aa",x"49",x"69"),
   887 => (x"7e",x"c1",x"87",x"c4"),
   888 => (x"ec",x"c0",x"87",x"d0"),
   889 => (x"87",x"c6",x"02",x"ad"),
   890 => (x"05",x"ad",x"fb",x"c0"),
   891 => (x"4b",x"c0",x"87",x"c4"),
   892 => (x"02",x"6e",x"7e",x"c1"),
   893 => (x"fa",x"87",x"f5",x"fe"),
   894 => (x"48",x"73",x"87",x"fd"),
   895 => (x"4d",x"26",x"8e",x"f8"),
   896 => (x"4b",x"26",x"4c",x"26"),
   897 => (x"00",x"00",x"4f",x"26"),
   898 => (x"1e",x"73",x"1e",x"00"),
   899 => (x"c8",x"4b",x"d4",x"ff"),
   900 => (x"d0",x"ff",x"4a",x"66"),
   901 => (x"78",x"c5",x"c8",x"48"),
   902 => (x"c1",x"48",x"d4",x"ff"),
   903 => (x"7b",x"11",x"78",x"d4"),
   904 => (x"f9",x"05",x"8a",x"c1"),
   905 => (x"48",x"d0",x"ff",x"87"),
   906 => (x"4b",x"26",x"78",x"c4"),
   907 => (x"5e",x"0e",x"4f",x"26"),
   908 => (x"0e",x"5d",x"5c",x"5b"),
   909 => (x"7e",x"71",x"86",x"f8"),
   910 => (x"e5",x"c2",x"1e",x"6e"),
   911 => (x"da",x"e9",x"49",x"d4"),
   912 => (x"70",x"86",x"c4",x"87"),
   913 => (x"e4",x"c4",x"02",x"98"),
   914 => (x"c8",x"e6",x"c1",x"87"),
   915 => (x"49",x"6e",x"4c",x"bf"),
   916 => (x"c8",x"87",x"d5",x"fc"),
   917 => (x"98",x"70",x"58",x"a6"),
   918 => (x"c4",x"87",x"c5",x"05"),
   919 => (x"78",x"c1",x"48",x"a6"),
   920 => (x"c5",x"48",x"d0",x"ff"),
   921 => (x"48",x"d4",x"ff",x"78"),
   922 => (x"c4",x"78",x"d5",x"c1"),
   923 => (x"89",x"c1",x"49",x"66"),
   924 => (x"e6",x"c1",x"31",x"c6"),
   925 => (x"4a",x"bf",x"97",x"c0"),
   926 => (x"ff",x"b0",x"71",x"48"),
   927 => (x"ff",x"78",x"08",x"d4"),
   928 => (x"78",x"c4",x"48",x"d0"),
   929 => (x"97",x"d0",x"e5",x"c2"),
   930 => (x"99",x"d0",x"49",x"bf"),
   931 => (x"c5",x"87",x"dd",x"02"),
   932 => (x"48",x"d4",x"ff",x"78"),
   933 => (x"c0",x"78",x"d6",x"c1"),
   934 => (x"48",x"d4",x"ff",x"4a"),
   935 => (x"c1",x"78",x"ff",x"c3"),
   936 => (x"aa",x"e0",x"c0",x"82"),
   937 => (x"ff",x"87",x"f2",x"04"),
   938 => (x"78",x"c4",x"48",x"d0"),
   939 => (x"c3",x"48",x"d4",x"ff"),
   940 => (x"d0",x"ff",x"78",x"ff"),
   941 => (x"ff",x"78",x"c5",x"48"),
   942 => (x"d3",x"c1",x"48",x"d4"),
   943 => (x"ff",x"78",x"c1",x"78"),
   944 => (x"78",x"c4",x"48",x"d0"),
   945 => (x"06",x"ac",x"b7",x"c0"),
   946 => (x"c2",x"87",x"cb",x"c2"),
   947 => (x"4b",x"bf",x"dc",x"e5"),
   948 => (x"73",x"7e",x"74",x"8c"),
   949 => (x"dd",x"c1",x"02",x"9b"),
   950 => (x"4d",x"c0",x"c8",x"87"),
   951 => (x"ab",x"b7",x"c0",x"8b"),
   952 => (x"c8",x"87",x"c6",x"03"),
   953 => (x"c0",x"4d",x"a3",x"c0"),
   954 => (x"d0",x"e5",x"c2",x"4b"),
   955 => (x"d0",x"49",x"bf",x"97"),
   956 => (x"87",x"cf",x"02",x"99"),
   957 => (x"e5",x"c2",x"1e",x"c0"),
   958 => (x"c7",x"eb",x"49",x"d4"),
   959 => (x"70",x"86",x"c4",x"87"),
   960 => (x"c2",x"87",x"d8",x"4c"),
   961 => (x"c2",x"1e",x"d4",x"d8"),
   962 => (x"ea",x"49",x"d4",x"e5"),
   963 => (x"4c",x"70",x"87",x"f6"),
   964 => (x"d8",x"c2",x"1e",x"75"),
   965 => (x"f0",x"fb",x"49",x"d4"),
   966 => (x"74",x"86",x"c8",x"87"),
   967 => (x"87",x"c5",x"05",x"9c"),
   968 => (x"ca",x"c1",x"48",x"c0"),
   969 => (x"c2",x"1e",x"c1",x"87"),
   970 => (x"e9",x"49",x"d4",x"e5"),
   971 => (x"86",x"c4",x"87",x"c7"),
   972 => (x"fe",x"05",x"9b",x"73"),
   973 => (x"4c",x"6e",x"87",x"e3"),
   974 => (x"06",x"ac",x"b7",x"c0"),
   975 => (x"e5",x"c2",x"87",x"d1"),
   976 => (x"78",x"c0",x"48",x"d4"),
   977 => (x"78",x"c0",x"80",x"d0"),
   978 => (x"e5",x"c2",x"80",x"f4"),
   979 => (x"c0",x"78",x"bf",x"e0"),
   980 => (x"fd",x"01",x"ac",x"b7"),
   981 => (x"d0",x"ff",x"87",x"f5"),
   982 => (x"ff",x"78",x"c5",x"48"),
   983 => (x"d3",x"c1",x"48",x"d4"),
   984 => (x"ff",x"78",x"c0",x"78"),
   985 => (x"78",x"c4",x"48",x"d0"),
   986 => (x"c2",x"c0",x"48",x"c1"),
   987 => (x"f8",x"48",x"c0",x"87"),
   988 => (x"26",x"4d",x"26",x"8e"),
   989 => (x"26",x"4b",x"26",x"4c"),
   990 => (x"5b",x"5e",x"0e",x"4f"),
   991 => (x"fc",x"0e",x"5d",x"5c"),
   992 => (x"c0",x"4d",x"71",x"86"),
   993 => (x"04",x"ad",x"4c",x"4b"),
   994 => (x"c0",x"87",x"e8",x"c0"),
   995 => (x"74",x"1e",x"e8",x"f5"),
   996 => (x"87",x"c4",x"02",x"9c"),
   997 => (x"87",x"c2",x"4a",x"c0"),
   998 => (x"49",x"72",x"4a",x"c1"),
   999 => (x"c4",x"87",x"fd",x"eb"),
  1000 => (x"c1",x"7e",x"70",x"86"),
  1001 => (x"c2",x"05",x"6e",x"83"),
  1002 => (x"c1",x"4b",x"75",x"87"),
  1003 => (x"06",x"ab",x"75",x"84"),
  1004 => (x"6e",x"87",x"d8",x"ff"),
  1005 => (x"26",x"8e",x"fc",x"48"),
  1006 => (x"26",x"4c",x"26",x"4d"),
  1007 => (x"1e",x"4f",x"26",x"4b"),
  1008 => (x"66",x"c4",x"4a",x"71"),
  1009 => (x"72",x"87",x"c5",x"05"),
  1010 => (x"87",x"e2",x"f9",x"49"),
  1011 => (x"5e",x"0e",x"4f",x"26"),
  1012 => (x"0e",x"5d",x"5c",x"5b"),
  1013 => (x"4c",x"71",x"86",x"fc"),
  1014 => (x"c2",x"91",x"de",x"49"),
  1015 => (x"71",x"4d",x"c0",x"e6"),
  1016 => (x"02",x"6d",x"97",x"85"),
  1017 => (x"c2",x"87",x"dc",x"c1"),
  1018 => (x"49",x"bf",x"f0",x"e5"),
  1019 => (x"fe",x"71",x"81",x"74"),
  1020 => (x"7e",x"70",x"87",x"c7"),
  1021 => (x"c0",x"02",x"98",x"48"),
  1022 => (x"e5",x"c2",x"87",x"f2"),
  1023 => (x"4a",x"70",x"4b",x"f4"),
  1024 => (x"c4",x"ff",x"49",x"cb"),
  1025 => (x"4b",x"74",x"87",x"dd"),
  1026 => (x"e6",x"c1",x"93",x"cc"),
  1027 => (x"83",x"c4",x"83",x"cc"),
  1028 => (x"7b",x"d0",x"c1",x"c1"),
  1029 => (x"c3",x"c1",x"49",x"74"),
  1030 => (x"7b",x"75",x"87",x"fa"),
  1031 => (x"97",x"c4",x"e6",x"c1"),
  1032 => (x"c2",x"1e",x"49",x"bf"),
  1033 => (x"fe",x"49",x"f4",x"e5"),
  1034 => (x"86",x"c4",x"87",x"d5"),
  1035 => (x"c3",x"c1",x"49",x"74"),
  1036 => (x"49",x"c0",x"87",x"e2"),
  1037 => (x"87",x"fd",x"c4",x"c1"),
  1038 => (x"48",x"cc",x"e5",x"c2"),
  1039 => (x"c0",x"49",x"50",x"c0"),
  1040 => (x"fc",x"87",x"e6",x"e2"),
  1041 => (x"26",x"4d",x"26",x"8e"),
  1042 => (x"26",x"4b",x"26",x"4c"),
  1043 => (x"00",x"00",x"00",x"4f"),
  1044 => (x"64",x"61",x"6f",x"4c"),
  1045 => (x"2e",x"67",x"6e",x"69"),
  1046 => (x"00",x"00",x"2e",x"2e"),
  1047 => (x"61",x"42",x"20",x"80"),
  1048 => (x"00",x"00",x"6b",x"63"),
  1049 => (x"64",x"61",x"6f",x"4c"),
  1050 => (x"20",x"2e",x"2a",x"20"),
  1051 => (x"00",x"00",x"00",x"00"),
  1052 => (x"00",x"00",x"20",x"3a"),
  1053 => (x"61",x"42",x"20",x"80"),
  1054 => (x"00",x"00",x"6b",x"63"),
  1055 => (x"78",x"45",x"20",x"80"),
  1056 => (x"00",x"00",x"74",x"69"),
  1057 => (x"49",x"20",x"44",x"53"),
  1058 => (x"2e",x"74",x"69",x"6e"),
  1059 => (x"00",x"00",x"00",x"2e"),
  1060 => (x"00",x"00",x"4b",x"4f"),
  1061 => (x"54",x"4f",x"4f",x"42"),
  1062 => (x"20",x"20",x"20",x"20"),
  1063 => (x"00",x"4d",x"4f",x"52"),
  1064 => (x"71",x"1e",x"73",x"1e"),
  1065 => (x"e5",x"c2",x"49",x"4b"),
  1066 => (x"71",x"81",x"bf",x"f0"),
  1067 => (x"70",x"87",x"ca",x"fb"),
  1068 => (x"c4",x"02",x"9a",x"4a"),
  1069 => (x"e9",x"e6",x"49",x"87"),
  1070 => (x"f0",x"e5",x"c2",x"87"),
  1071 => (x"73",x"78",x"c0",x"48"),
  1072 => (x"87",x"fa",x"c1",x"49"),
  1073 => (x"4f",x"26",x"4b",x"26"),
  1074 => (x"71",x"1e",x"73",x"1e"),
  1075 => (x"4a",x"a3",x"c4",x"4b"),
  1076 => (x"87",x"d0",x"c1",x"02"),
  1077 => (x"dc",x"02",x"8a",x"c1"),
  1078 => (x"c0",x"02",x"8a",x"87"),
  1079 => (x"05",x"8a",x"87",x"f2"),
  1080 => (x"c2",x"87",x"d3",x"c1"),
  1081 => (x"02",x"bf",x"f0",x"e5"),
  1082 => (x"48",x"87",x"cb",x"c1"),
  1083 => (x"e5",x"c2",x"88",x"c1"),
  1084 => (x"c1",x"c1",x"58",x"f4"),
  1085 => (x"f0",x"e5",x"c2",x"87"),
  1086 => (x"89",x"c6",x"49",x"bf"),
  1087 => (x"59",x"f4",x"e5",x"c2"),
  1088 => (x"03",x"a9",x"b7",x"c0"),
  1089 => (x"c2",x"87",x"ef",x"c0"),
  1090 => (x"c0",x"48",x"f0",x"e5"),
  1091 => (x"87",x"e6",x"c0",x"78"),
  1092 => (x"bf",x"ec",x"e5",x"c2"),
  1093 => (x"c2",x"87",x"df",x"02"),
  1094 => (x"48",x"bf",x"f0",x"e5"),
  1095 => (x"e5",x"c2",x"80",x"c1"),
  1096 => (x"87",x"d2",x"58",x"f4"),
  1097 => (x"bf",x"ec",x"e5",x"c2"),
  1098 => (x"c2",x"87",x"cb",x"02"),
  1099 => (x"48",x"bf",x"f0",x"e5"),
  1100 => (x"e5",x"c2",x"80",x"c6"),
  1101 => (x"49",x"73",x"58",x"f4"),
  1102 => (x"4b",x"26",x"87",x"c4"),
  1103 => (x"5e",x"0e",x"4f",x"26"),
  1104 => (x"0e",x"5d",x"5c",x"5b"),
  1105 => (x"a6",x"d0",x"86",x"f0"),
  1106 => (x"d4",x"d8",x"c2",x"59"),
  1107 => (x"c2",x"4c",x"c0",x"4d"),
  1108 => (x"c1",x"48",x"ec",x"e5"),
  1109 => (x"48",x"a6",x"c8",x"78"),
  1110 => (x"7e",x"75",x"78",x"c0"),
  1111 => (x"bf",x"f0",x"e5",x"c2"),
  1112 => (x"06",x"a8",x"c0",x"48"),
  1113 => (x"c8",x"87",x"c0",x"c1"),
  1114 => (x"7e",x"75",x"5c",x"a6"),
  1115 => (x"48",x"d4",x"d8",x"c2"),
  1116 => (x"f2",x"c0",x"02",x"98"),
  1117 => (x"4d",x"66",x"c4",x"87"),
  1118 => (x"1e",x"e8",x"f5",x"c0"),
  1119 => (x"c4",x"02",x"66",x"cc"),
  1120 => (x"c2",x"4c",x"c0",x"87"),
  1121 => (x"74",x"4c",x"c1",x"87"),
  1122 => (x"87",x"d0",x"e4",x"49"),
  1123 => (x"7e",x"70",x"86",x"c4"),
  1124 => (x"66",x"c8",x"85",x"c1"),
  1125 => (x"cc",x"80",x"c1",x"48"),
  1126 => (x"e5",x"c2",x"58",x"a6"),
  1127 => (x"03",x"ad",x"bf",x"f0"),
  1128 => (x"05",x"6e",x"87",x"c5"),
  1129 => (x"6e",x"87",x"d1",x"ff"),
  1130 => (x"75",x"4c",x"c0",x"4d"),
  1131 => (x"dc",x"c3",x"02",x"9d"),
  1132 => (x"e8",x"f5",x"c0",x"87"),
  1133 => (x"02",x"66",x"cc",x"1e"),
  1134 => (x"a6",x"c8",x"87",x"c7"),
  1135 => (x"c5",x"78",x"c0",x"48"),
  1136 => (x"48",x"a6",x"c8",x"87"),
  1137 => (x"66",x"c8",x"78",x"c1"),
  1138 => (x"87",x"d0",x"e3",x"49"),
  1139 => (x"7e",x"70",x"86",x"c4"),
  1140 => (x"c2",x"02",x"98",x"48"),
  1141 => (x"cb",x"49",x"87",x"e4"),
  1142 => (x"49",x"69",x"97",x"81"),
  1143 => (x"c1",x"02",x"99",x"d0"),
  1144 => (x"49",x"74",x"87",x"d4"),
  1145 => (x"e6",x"c1",x"91",x"cc"),
  1146 => (x"c2",x"c1",x"81",x"cc"),
  1147 => (x"81",x"c8",x"79",x"e0"),
  1148 => (x"74",x"51",x"ff",x"c3"),
  1149 => (x"c2",x"91",x"de",x"49"),
  1150 => (x"71",x"4d",x"c0",x"e6"),
  1151 => (x"97",x"c1",x"c2",x"85"),
  1152 => (x"49",x"a5",x"c1",x"7d"),
  1153 => (x"c2",x"51",x"e0",x"c0"),
  1154 => (x"bf",x"97",x"e4",x"e0"),
  1155 => (x"c1",x"87",x"d2",x"02"),
  1156 => (x"4b",x"a5",x"c2",x"84"),
  1157 => (x"4a",x"e4",x"e0",x"c2"),
  1158 => (x"fc",x"fe",x"49",x"db"),
  1159 => (x"d9",x"c1",x"87",x"c5"),
  1160 => (x"49",x"a5",x"cd",x"87"),
  1161 => (x"84",x"c1",x"51",x"c0"),
  1162 => (x"6e",x"4b",x"a5",x"c2"),
  1163 => (x"fe",x"49",x"cb",x"4a"),
  1164 => (x"c1",x"87",x"f0",x"fb"),
  1165 => (x"49",x"74",x"87",x"c4"),
  1166 => (x"e6",x"c1",x"91",x"cc"),
  1167 => (x"ff",x"c0",x"81",x"cc"),
  1168 => (x"e0",x"c2",x"79",x"ce"),
  1169 => (x"02",x"bf",x"97",x"e4"),
  1170 => (x"49",x"74",x"87",x"d8"),
  1171 => (x"84",x"c1",x"91",x"de"),
  1172 => (x"4b",x"c0",x"e6",x"c2"),
  1173 => (x"e0",x"c2",x"83",x"71"),
  1174 => (x"49",x"dd",x"4a",x"e4"),
  1175 => (x"87",x"c3",x"fb",x"fe"),
  1176 => (x"4b",x"74",x"87",x"d8"),
  1177 => (x"e6",x"c2",x"93",x"de"),
  1178 => (x"a3",x"cb",x"83",x"c0"),
  1179 => (x"c1",x"51",x"c0",x"49"),
  1180 => (x"4a",x"6e",x"73",x"84"),
  1181 => (x"fa",x"fe",x"49",x"cb"),
  1182 => (x"66",x"c8",x"87",x"e9"),
  1183 => (x"cc",x"80",x"c1",x"48"),
  1184 => (x"ac",x"c7",x"58",x"a6"),
  1185 => (x"87",x"c5",x"c0",x"03"),
  1186 => (x"e4",x"fc",x"05",x"6e"),
  1187 => (x"03",x"ac",x"c7",x"87"),
  1188 => (x"c2",x"87",x"e4",x"c0"),
  1189 => (x"c0",x"48",x"ec",x"e5"),
  1190 => (x"cc",x"49",x"74",x"78"),
  1191 => (x"cc",x"e6",x"c1",x"91"),
  1192 => (x"ce",x"ff",x"c0",x"81"),
  1193 => (x"de",x"49",x"74",x"79"),
  1194 => (x"c0",x"e6",x"c2",x"91"),
  1195 => (x"c1",x"51",x"c0",x"81"),
  1196 => (x"04",x"ac",x"c7",x"84"),
  1197 => (x"c1",x"87",x"dc",x"ff"),
  1198 => (x"c0",x"48",x"e8",x"e7"),
  1199 => (x"c1",x"80",x"f7",x"50"),
  1200 => (x"c1",x"40",x"e4",x"cc"),
  1201 => (x"c8",x"78",x"dc",x"c1"),
  1202 => (x"c8",x"c3",x"c1",x"80"),
  1203 => (x"49",x"66",x"cc",x"78"),
  1204 => (x"87",x"c0",x"f9",x"c0"),
  1205 => (x"4d",x"26",x"8e",x"f0"),
  1206 => (x"4b",x"26",x"4c",x"26"),
  1207 => (x"73",x"1e",x"4f",x"26"),
  1208 => (x"49",x"4b",x"71",x"1e"),
  1209 => (x"e6",x"c1",x"91",x"cc"),
  1210 => (x"a1",x"c8",x"81",x"cc"),
  1211 => (x"c0",x"e6",x"c1",x"4a"),
  1212 => (x"c9",x"50",x"12",x"48"),
  1213 => (x"f8",x"c0",x"4a",x"a1"),
  1214 => (x"50",x"12",x"48",x"c8"),
  1215 => (x"e6",x"c1",x"81",x"ca"),
  1216 => (x"50",x"11",x"48",x"c4"),
  1217 => (x"97",x"c4",x"e6",x"c1"),
  1218 => (x"c0",x"1e",x"49",x"bf"),
  1219 => (x"87",x"ef",x"f2",x"49"),
  1220 => (x"e9",x"f8",x"49",x"73"),
  1221 => (x"26",x"8e",x"fc",x"87"),
  1222 => (x"1e",x"4f",x"26",x"4b"),
  1223 => (x"f9",x"c0",x"49",x"c0"),
  1224 => (x"4f",x"26",x"87",x"d3"),
  1225 => (x"49",x"4a",x"71",x"1e"),
  1226 => (x"e6",x"c1",x"91",x"cc"),
  1227 => (x"81",x"c8",x"81",x"cc"),
  1228 => (x"48",x"cc",x"e5",x"c2"),
  1229 => (x"f0",x"c0",x"50",x"11"),
  1230 => (x"f5",x"fe",x"49",x"a2"),
  1231 => (x"49",x"c0",x"87",x"ce"),
  1232 => (x"26",x"87",x"e6",x"d6"),
  1233 => (x"d4",x"ff",x"1e",x"4f"),
  1234 => (x"7a",x"ff",x"c3",x"4a"),
  1235 => (x"c0",x"48",x"d0",x"ff"),
  1236 => (x"7a",x"de",x"78",x"e1"),
  1237 => (x"c8",x"48",x"7a",x"71"),
  1238 => (x"7a",x"70",x"28",x"b7"),
  1239 => (x"b7",x"d0",x"48",x"71"),
  1240 => (x"71",x"7a",x"70",x"28"),
  1241 => (x"28",x"b7",x"d8",x"48"),
  1242 => (x"d0",x"ff",x"7a",x"70"),
  1243 => (x"78",x"e0",x"c0",x"48"),
  1244 => (x"5e",x"0e",x"4f",x"26"),
  1245 => (x"0e",x"5d",x"5c",x"5b"),
  1246 => (x"4d",x"71",x"86",x"f4"),
  1247 => (x"c1",x"91",x"cc",x"49"),
  1248 => (x"c8",x"81",x"cc",x"e6"),
  1249 => (x"a1",x"ca",x"4a",x"a1"),
  1250 => (x"48",x"a6",x"c4",x"7e"),
  1251 => (x"bf",x"c8",x"e5",x"c2"),
  1252 => (x"bf",x"97",x"6e",x"78"),
  1253 => (x"4c",x"66",x"c4",x"4b"),
  1254 => (x"48",x"12",x"2c",x"73"),
  1255 => (x"70",x"58",x"a6",x"cc"),
  1256 => (x"c9",x"84",x"c1",x"9c"),
  1257 => (x"49",x"69",x"97",x"81"),
  1258 => (x"c2",x"04",x"ac",x"b7"),
  1259 => (x"6e",x"4c",x"c0",x"87"),
  1260 => (x"c8",x"4a",x"bf",x"97"),
  1261 => (x"31",x"72",x"49",x"66"),
  1262 => (x"66",x"c4",x"b9",x"ff"),
  1263 => (x"72",x"48",x"74",x"99"),
  1264 => (x"b1",x"4a",x"70",x"30"),
  1265 => (x"59",x"cc",x"e5",x"c2"),
  1266 => (x"87",x"f9",x"fd",x"71"),
  1267 => (x"e5",x"c2",x"1e",x"c7"),
  1268 => (x"c1",x"1e",x"bf",x"e8"),
  1269 => (x"c2",x"1e",x"cc",x"e6"),
  1270 => (x"bf",x"97",x"cc",x"e5"),
  1271 => (x"87",x"f4",x"c1",x"49"),
  1272 => (x"f4",x"c0",x"49",x"75"),
  1273 => (x"8e",x"e8",x"87",x"ee"),
  1274 => (x"4c",x"26",x"4d",x"26"),
  1275 => (x"4f",x"26",x"4b",x"26"),
  1276 => (x"71",x"1e",x"73",x"1e"),
  1277 => (x"f9",x"fd",x"49",x"4b"),
  1278 => (x"fd",x"49",x"73",x"87"),
  1279 => (x"4b",x"26",x"87",x"f4"),
  1280 => (x"73",x"1e",x"4f",x"26"),
  1281 => (x"c2",x"4b",x"71",x"1e"),
  1282 => (x"d6",x"02",x"4a",x"a3"),
  1283 => (x"05",x"8a",x"c1",x"87"),
  1284 => (x"c2",x"87",x"e2",x"c0"),
  1285 => (x"02",x"bf",x"e8",x"e5"),
  1286 => (x"c1",x"48",x"87",x"db"),
  1287 => (x"ec",x"e5",x"c2",x"88"),
  1288 => (x"c2",x"87",x"d2",x"58"),
  1289 => (x"02",x"bf",x"ec",x"e5"),
  1290 => (x"e5",x"c2",x"87",x"cb"),
  1291 => (x"c1",x"48",x"bf",x"e8"),
  1292 => (x"ec",x"e5",x"c2",x"80"),
  1293 => (x"c2",x"1e",x"c7",x"58"),
  1294 => (x"1e",x"bf",x"e8",x"e5"),
  1295 => (x"1e",x"cc",x"e6",x"c1"),
  1296 => (x"97",x"cc",x"e5",x"c2"),
  1297 => (x"87",x"cc",x"49",x"bf"),
  1298 => (x"f3",x"c0",x"49",x"73"),
  1299 => (x"8e",x"f4",x"87",x"c6"),
  1300 => (x"4f",x"26",x"4b",x"26"),
  1301 => (x"5c",x"5b",x"5e",x"0e"),
  1302 => (x"cc",x"ff",x"0e",x"5d"),
  1303 => (x"a6",x"e4",x"c0",x"86"),
  1304 => (x"48",x"a6",x"cc",x"59"),
  1305 => (x"80",x"c4",x"78",x"c0"),
  1306 => (x"80",x"c4",x"78",x"c0"),
  1307 => (x"78",x"66",x"c8",x"c1"),
  1308 => (x"78",x"c1",x"80",x"c4"),
  1309 => (x"78",x"c1",x"80",x"c4"),
  1310 => (x"48",x"ec",x"e5",x"c2"),
  1311 => (x"e2",x"e0",x"78",x"c1"),
  1312 => (x"87",x"fc",x"e0",x"87"),
  1313 => (x"70",x"87",x"d1",x"e0"),
  1314 => (x"ac",x"fb",x"c0",x"4c"),
  1315 => (x"87",x"f3",x"c1",x"02"),
  1316 => (x"05",x"66",x"e0",x"c0"),
  1317 => (x"c1",x"87",x"e8",x"c1"),
  1318 => (x"c4",x"4a",x"66",x"c4"),
  1319 => (x"c1",x"7e",x"6a",x"82"),
  1320 => (x"6e",x"48",x"e4",x"c1"),
  1321 => (x"20",x"41",x"20",x"49"),
  1322 => (x"c1",x"51",x"10",x"41"),
  1323 => (x"c1",x"48",x"66",x"c4"),
  1324 => (x"6a",x"78",x"de",x"cb"),
  1325 => (x"74",x"81",x"c7",x"49"),
  1326 => (x"66",x"c4",x"c1",x"51"),
  1327 => (x"c1",x"81",x"c8",x"49"),
  1328 => (x"48",x"a6",x"d8",x"51"),
  1329 => (x"c4",x"c1",x"78",x"c2"),
  1330 => (x"81",x"c9",x"49",x"66"),
  1331 => (x"c4",x"c1",x"51",x"c0"),
  1332 => (x"81",x"ca",x"49",x"66"),
  1333 => (x"1e",x"c1",x"51",x"c0"),
  1334 => (x"49",x"6a",x"1e",x"d8"),
  1335 => (x"df",x"ff",x"81",x"c8"),
  1336 => (x"86",x"c8",x"87",x"f2"),
  1337 => (x"48",x"66",x"c8",x"c1"),
  1338 => (x"c7",x"01",x"a8",x"c0"),
  1339 => (x"48",x"a6",x"d0",x"87"),
  1340 => (x"87",x"cf",x"78",x"c1"),
  1341 => (x"48",x"66",x"c8",x"c1"),
  1342 => (x"a6",x"d8",x"88",x"c1"),
  1343 => (x"ff",x"87",x"c4",x"58"),
  1344 => (x"74",x"87",x"fd",x"de"),
  1345 => (x"da",x"cd",x"02",x"9c"),
  1346 => (x"48",x"66",x"d0",x"87"),
  1347 => (x"a8",x"66",x"cc",x"c1"),
  1348 => (x"87",x"cf",x"cd",x"03"),
  1349 => (x"c0",x"48",x"a6",x"c8"),
  1350 => (x"dd",x"ff",x"7e",x"78"),
  1351 => (x"4c",x"70",x"87",x"fa"),
  1352 => (x"05",x"ac",x"d0",x"c1"),
  1353 => (x"c4",x"87",x"e7",x"c2"),
  1354 => (x"78",x"6e",x"48",x"a6"),
  1355 => (x"70",x"87",x"d0",x"e0"),
  1356 => (x"66",x"cc",x"48",x"7e"),
  1357 => (x"87",x"c5",x"06",x"a8"),
  1358 => (x"6e",x"48",x"a6",x"cc"),
  1359 => (x"d7",x"dd",x"ff",x"78"),
  1360 => (x"c0",x"4c",x"70",x"87"),
  1361 => (x"c1",x"05",x"ac",x"ec"),
  1362 => (x"66",x"d0",x"87",x"ee"),
  1363 => (x"c1",x"91",x"cc",x"49"),
  1364 => (x"c4",x"81",x"66",x"c4"),
  1365 => (x"4d",x"6a",x"4a",x"a1"),
  1366 => (x"6e",x"4a",x"a1",x"c8"),
  1367 => (x"e4",x"cc",x"c1",x"52"),
  1368 => (x"f3",x"dc",x"ff",x"79"),
  1369 => (x"9c",x"4c",x"70",x"87"),
  1370 => (x"c0",x"87",x"d9",x"02"),
  1371 => (x"d3",x"02",x"ac",x"fb"),
  1372 => (x"ff",x"55",x"74",x"87"),
  1373 => (x"70",x"87",x"e1",x"dc"),
  1374 => (x"c7",x"02",x"9c",x"4c"),
  1375 => (x"ac",x"fb",x"c0",x"87"),
  1376 => (x"87",x"ed",x"ff",x"05"),
  1377 => (x"c2",x"55",x"e0",x"c0"),
  1378 => (x"97",x"c0",x"55",x"c1"),
  1379 => (x"66",x"e0",x"c0",x"7d"),
  1380 => (x"a8",x"66",x"c4",x"48"),
  1381 => (x"d0",x"87",x"db",x"05"),
  1382 => (x"66",x"d4",x"48",x"66"),
  1383 => (x"87",x"ca",x"04",x"a8"),
  1384 => (x"c1",x"48",x"66",x"d0"),
  1385 => (x"58",x"a6",x"d4",x"80"),
  1386 => (x"66",x"d4",x"87",x"c8"),
  1387 => (x"d8",x"88",x"c1",x"48"),
  1388 => (x"db",x"ff",x"58",x"a6"),
  1389 => (x"4c",x"70",x"87",x"e2"),
  1390 => (x"05",x"ac",x"d0",x"c1"),
  1391 => (x"66",x"dc",x"87",x"c9"),
  1392 => (x"c0",x"80",x"c1",x"48"),
  1393 => (x"c1",x"58",x"a6",x"e0"),
  1394 => (x"fd",x"02",x"ac",x"d0"),
  1395 => (x"48",x"6e",x"87",x"d9"),
  1396 => (x"a8",x"66",x"e0",x"c0"),
  1397 => (x"87",x"eb",x"c9",x"05"),
  1398 => (x"48",x"a6",x"e4",x"c0"),
  1399 => (x"48",x"74",x"78",x"c0"),
  1400 => (x"c8",x"88",x"fb",x"c0"),
  1401 => (x"98",x"70",x"58",x"a6"),
  1402 => (x"87",x"dd",x"c9",x"02"),
  1403 => (x"c8",x"88",x"cb",x"48"),
  1404 => (x"98",x"70",x"58",x"a6"),
  1405 => (x"87",x"cf",x"c1",x"02"),
  1406 => (x"c8",x"88",x"c9",x"48"),
  1407 => (x"98",x"70",x"58",x"a6"),
  1408 => (x"87",x"ff",x"c3",x"02"),
  1409 => (x"c8",x"88",x"c4",x"48"),
  1410 => (x"98",x"70",x"58",x"a6"),
  1411 => (x"48",x"87",x"cf",x"02"),
  1412 => (x"a6",x"c8",x"88",x"c1"),
  1413 => (x"02",x"98",x"70",x"58"),
  1414 => (x"c8",x"87",x"e8",x"c3"),
  1415 => (x"a6",x"c8",x"87",x"dc"),
  1416 => (x"78",x"f0",x"c0",x"48"),
  1417 => (x"87",x"f0",x"d9",x"ff"),
  1418 => (x"ec",x"c0",x"4c",x"70"),
  1419 => (x"c3",x"c0",x"02",x"ac"),
  1420 => (x"5c",x"a6",x"cc",x"87"),
  1421 => (x"02",x"ac",x"ec",x"c0"),
  1422 => (x"d9",x"ff",x"87",x"cd"),
  1423 => (x"4c",x"70",x"87",x"da"),
  1424 => (x"05",x"ac",x"ec",x"c0"),
  1425 => (x"c0",x"87",x"f3",x"ff"),
  1426 => (x"c0",x"02",x"ac",x"ec"),
  1427 => (x"d9",x"ff",x"87",x"c4"),
  1428 => (x"1e",x"c0",x"87",x"c6"),
  1429 => (x"66",x"d8",x"1e",x"ca"),
  1430 => (x"c1",x"91",x"cc",x"49"),
  1431 => (x"71",x"48",x"66",x"cc"),
  1432 => (x"58",x"a6",x"cc",x"80"),
  1433 => (x"c4",x"48",x"66",x"c8"),
  1434 => (x"58",x"a6",x"d0",x"80"),
  1435 => (x"49",x"bf",x"66",x"cc"),
  1436 => (x"87",x"e0",x"d9",x"ff"),
  1437 => (x"1e",x"de",x"1e",x"c1"),
  1438 => (x"49",x"bf",x"66",x"d4"),
  1439 => (x"87",x"d4",x"d9",x"ff"),
  1440 => (x"49",x"70",x"86",x"d0"),
  1441 => (x"88",x"08",x"c0",x"48"),
  1442 => (x"58",x"a6",x"ec",x"c0"),
  1443 => (x"c0",x"06",x"a8",x"c0"),
  1444 => (x"e8",x"c0",x"87",x"ee"),
  1445 => (x"a8",x"dd",x"48",x"66"),
  1446 => (x"87",x"e4",x"c0",x"03"),
  1447 => (x"49",x"bf",x"66",x"c4"),
  1448 => (x"81",x"66",x"e8",x"c0"),
  1449 => (x"c0",x"51",x"e0",x"c0"),
  1450 => (x"c1",x"49",x"66",x"e8"),
  1451 => (x"bf",x"66",x"c4",x"81"),
  1452 => (x"51",x"c1",x"c2",x"81"),
  1453 => (x"49",x"66",x"e8",x"c0"),
  1454 => (x"66",x"c4",x"81",x"c2"),
  1455 => (x"51",x"c0",x"81",x"bf"),
  1456 => (x"cb",x"c1",x"48",x"6e"),
  1457 => (x"49",x"6e",x"78",x"de"),
  1458 => (x"66",x"d8",x"81",x"c8"),
  1459 => (x"c9",x"49",x"6e",x"51"),
  1460 => (x"51",x"66",x"dc",x"81"),
  1461 => (x"81",x"ca",x"49",x"6e"),
  1462 => (x"d8",x"51",x"66",x"c8"),
  1463 => (x"80",x"c1",x"48",x"66"),
  1464 => (x"d0",x"58",x"a6",x"dc"),
  1465 => (x"66",x"d4",x"48",x"66"),
  1466 => (x"cb",x"c0",x"04",x"a8"),
  1467 => (x"48",x"66",x"d0",x"87"),
  1468 => (x"a6",x"d4",x"80",x"c1"),
  1469 => (x"87",x"d1",x"c5",x"58"),
  1470 => (x"c1",x"48",x"66",x"d4"),
  1471 => (x"58",x"a6",x"d8",x"88"),
  1472 => (x"ff",x"87",x"c6",x"c5"),
  1473 => (x"c0",x"87",x"f8",x"d8"),
  1474 => (x"ff",x"58",x"a6",x"ec"),
  1475 => (x"c0",x"87",x"f0",x"d8"),
  1476 => (x"c0",x"58",x"a6",x"f0"),
  1477 => (x"c0",x"05",x"a8",x"ec"),
  1478 => (x"48",x"a6",x"87",x"c9"),
  1479 => (x"78",x"66",x"e8",x"c0"),
  1480 => (x"ff",x"87",x"c4",x"c0"),
  1481 => (x"d0",x"87",x"f1",x"d5"),
  1482 => (x"91",x"cc",x"49",x"66"),
  1483 => (x"48",x"66",x"c4",x"c1"),
  1484 => (x"a6",x"c8",x"80",x"71"),
  1485 => (x"4a",x"66",x"c4",x"58"),
  1486 => (x"66",x"c4",x"82",x"c8"),
  1487 => (x"c0",x"81",x"ca",x"49"),
  1488 => (x"c0",x"51",x"66",x"e8"),
  1489 => (x"c1",x"49",x"66",x"ec"),
  1490 => (x"66",x"e8",x"c0",x"81"),
  1491 => (x"71",x"48",x"c1",x"89"),
  1492 => (x"c1",x"49",x"70",x"30"),
  1493 => (x"7a",x"97",x"71",x"89"),
  1494 => (x"bf",x"c8",x"e5",x"c2"),
  1495 => (x"66",x"e8",x"c0",x"49"),
  1496 => (x"4a",x"6a",x"97",x"29"),
  1497 => (x"c0",x"98",x"71",x"48"),
  1498 => (x"c4",x"58",x"a6",x"f4"),
  1499 => (x"80",x"c4",x"48",x"66"),
  1500 => (x"c8",x"58",x"a6",x"cc"),
  1501 => (x"c0",x"4d",x"bf",x"66"),
  1502 => (x"6e",x"48",x"66",x"e0"),
  1503 => (x"c5",x"c0",x"02",x"a8"),
  1504 => (x"c0",x"7e",x"c0",x"87"),
  1505 => (x"7e",x"c1",x"87",x"c2"),
  1506 => (x"e0",x"c0",x"1e",x"6e"),
  1507 => (x"ff",x"49",x"75",x"1e"),
  1508 => (x"c8",x"87",x"c1",x"d5"),
  1509 => (x"c0",x"4c",x"70",x"86"),
  1510 => (x"c1",x"06",x"ac",x"b7"),
  1511 => (x"85",x"74",x"87",x"d4"),
  1512 => (x"49",x"bf",x"66",x"c8"),
  1513 => (x"75",x"81",x"e0",x"c0"),
  1514 => (x"c1",x"c1",x"4b",x"89"),
  1515 => (x"fe",x"71",x"4a",x"f0"),
  1516 => (x"c2",x"87",x"f0",x"e5"),
  1517 => (x"c0",x"7e",x"75",x"85"),
  1518 => (x"c1",x"48",x"66",x"e4"),
  1519 => (x"a6",x"e8",x"c0",x"80"),
  1520 => (x"66",x"f0",x"c0",x"58"),
  1521 => (x"70",x"81",x"c1",x"49"),
  1522 => (x"c5",x"c0",x"02",x"a9"),
  1523 => (x"c0",x"4d",x"c0",x"87"),
  1524 => (x"4d",x"c1",x"87",x"c2"),
  1525 => (x"66",x"cc",x"1e",x"75"),
  1526 => (x"e0",x"c0",x"49",x"bf"),
  1527 => (x"89",x"66",x"c4",x"81"),
  1528 => (x"66",x"c8",x"1e",x"71"),
  1529 => (x"eb",x"d3",x"ff",x"49"),
  1530 => (x"c0",x"86",x"c8",x"87"),
  1531 => (x"ff",x"01",x"a8",x"b7"),
  1532 => (x"e4",x"c0",x"87",x"c5"),
  1533 => (x"d3",x"c0",x"02",x"66"),
  1534 => (x"49",x"66",x"c4",x"87"),
  1535 => (x"e4",x"c0",x"81",x"c9"),
  1536 => (x"66",x"c4",x"51",x"66"),
  1537 => (x"f2",x"cd",x"c1",x"48"),
  1538 => (x"87",x"ce",x"c0",x"78"),
  1539 => (x"c9",x"49",x"66",x"c4"),
  1540 => (x"c4",x"51",x"c2",x"81"),
  1541 => (x"cf",x"c1",x"48",x"66"),
  1542 => (x"66",x"d0",x"78",x"f0"),
  1543 => (x"a8",x"66",x"d4",x"48"),
  1544 => (x"87",x"cb",x"c0",x"04"),
  1545 => (x"c1",x"48",x"66",x"d0"),
  1546 => (x"58",x"a6",x"d4",x"80"),
  1547 => (x"d4",x"87",x"da",x"c0"),
  1548 => (x"88",x"c1",x"48",x"66"),
  1549 => (x"c0",x"58",x"a6",x"d8"),
  1550 => (x"d2",x"ff",x"87",x"cf"),
  1551 => (x"4c",x"70",x"87",x"c2"),
  1552 => (x"ff",x"87",x"c6",x"c0"),
  1553 => (x"70",x"87",x"f9",x"d1"),
  1554 => (x"48",x"66",x"dc",x"4c"),
  1555 => (x"e0",x"c0",x"80",x"c1"),
  1556 => (x"9c",x"74",x"58",x"a6"),
  1557 => (x"87",x"cb",x"c0",x"02"),
  1558 => (x"c1",x"48",x"66",x"d0"),
  1559 => (x"04",x"a8",x"66",x"cc"),
  1560 => (x"d0",x"87",x"f1",x"f2"),
  1561 => (x"a8",x"c7",x"48",x"66"),
  1562 => (x"87",x"e1",x"c0",x"03"),
  1563 => (x"c2",x"4c",x"66",x"d0"),
  1564 => (x"c0",x"48",x"ec",x"e5"),
  1565 => (x"cc",x"49",x"74",x"78"),
  1566 => (x"66",x"c4",x"c1",x"91"),
  1567 => (x"4a",x"a1",x"c4",x"81"),
  1568 => (x"52",x"c0",x"4a",x"6a"),
  1569 => (x"c7",x"84",x"c1",x"79"),
  1570 => (x"e2",x"ff",x"04",x"ac"),
  1571 => (x"66",x"e0",x"c0",x"87"),
  1572 => (x"87",x"e2",x"c0",x"02"),
  1573 => (x"49",x"66",x"c4",x"c1"),
  1574 => (x"c1",x"81",x"d4",x"c1"),
  1575 => (x"c1",x"4a",x"66",x"c4"),
  1576 => (x"52",x"c0",x"82",x"dc"),
  1577 => (x"79",x"e4",x"cc",x"c1"),
  1578 => (x"49",x"66",x"c4",x"c1"),
  1579 => (x"c1",x"81",x"d8",x"c1"),
  1580 => (x"c0",x"79",x"f4",x"c1"),
  1581 => (x"c4",x"c1",x"87",x"d6"),
  1582 => (x"d4",x"c1",x"49",x"66"),
  1583 => (x"66",x"c4",x"c1",x"81"),
  1584 => (x"82",x"d8",x"c1",x"4a"),
  1585 => (x"7a",x"fc",x"c1",x"c1"),
  1586 => (x"79",x"db",x"cc",x"c1"),
  1587 => (x"49",x"66",x"c4",x"c1"),
  1588 => (x"c1",x"81",x"e0",x"c1"),
  1589 => (x"ff",x"79",x"c2",x"d0"),
  1590 => (x"cc",x"87",x"dc",x"cf"),
  1591 => (x"cc",x"ff",x"48",x"66"),
  1592 => (x"26",x"4d",x"26",x"8e"),
  1593 => (x"26",x"4b",x"26",x"4c"),
  1594 => (x"1e",x"c7",x"1e",x"4f"),
  1595 => (x"bf",x"e8",x"e5",x"c2"),
  1596 => (x"cc",x"e6",x"c1",x"1e"),
  1597 => (x"cc",x"e5",x"c2",x"1e"),
  1598 => (x"ed",x"49",x"bf",x"97"),
  1599 => (x"e6",x"c1",x"87",x"d6"),
  1600 => (x"e1",x"c0",x"49",x"cc"),
  1601 => (x"8e",x"f4",x"87",x"dc"),
  1602 => (x"73",x"1e",x"4f",x"26"),
  1603 => (x"87",x"d9",x"c7",x"1e"),
  1604 => (x"48",x"f4",x"e5",x"c2"),
  1605 => (x"d4",x"ff",x"50",x"c0"),
  1606 => (x"78",x"ff",x"c3",x"48"),
  1607 => (x"49",x"c4",x"c2",x"c1"),
  1608 => (x"87",x"c3",x"de",x"fe"),
  1609 => (x"87",x"d8",x"e9",x"fe"),
  1610 => (x"cd",x"02",x"98",x"70"),
  1611 => (x"cb",x"f1",x"fe",x"87"),
  1612 => (x"02",x"98",x"70",x"87"),
  1613 => (x"4a",x"c1",x"87",x"c4"),
  1614 => (x"4a",x"c0",x"87",x"c2"),
  1615 => (x"c8",x"02",x"9a",x"72"),
  1616 => (x"d0",x"c2",x"c1",x"87"),
  1617 => (x"de",x"dd",x"fe",x"49"),
  1618 => (x"e8",x"e5",x"c2",x"87"),
  1619 => (x"c2",x"78",x"c0",x"48"),
  1620 => (x"c0",x"48",x"cc",x"e5"),
  1621 => (x"d0",x"fe",x"49",x"50"),
  1622 => (x"fc",x"ef",x"c0",x"87"),
  1623 => (x"9b",x"4b",x"70",x"87"),
  1624 => (x"c1",x"87",x"cf",x"02"),
  1625 => (x"c7",x"5b",x"e8",x"e7"),
  1626 => (x"87",x"e8",x"de",x"49"),
  1627 => (x"e0",x"c0",x"49",x"c1"),
  1628 => (x"ee",x"c2",x"87",x"c3"),
  1629 => (x"e4",x"e1",x"c0",x"87"),
  1630 => (x"26",x"87",x"fa",x"87"),
  1631 => (x"00",x"4f",x"26",x"4b"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"00",x"01"),
  1635 => (x"00",x"00",x"0f",x"ce"),
  1636 => (x"00",x"00",x"29",x"80"),
  1637 => (x"00",x"00",x"00",x"00"),
  1638 => (x"00",x"00",x"0f",x"ce"),
  1639 => (x"00",x"00",x"29",x"9e"),
  1640 => (x"00",x"00",x"00",x"00"),
  1641 => (x"00",x"00",x"0f",x"ce"),
  1642 => (x"00",x"00",x"29",x"bc"),
  1643 => (x"00",x"00",x"00",x"00"),
  1644 => (x"00",x"00",x"0f",x"ce"),
  1645 => (x"00",x"00",x"29",x"da"),
  1646 => (x"00",x"00",x"00",x"00"),
  1647 => (x"00",x"00",x"0f",x"ce"),
  1648 => (x"00",x"00",x"29",x"f8"),
  1649 => (x"00",x"00",x"00",x"00"),
  1650 => (x"00",x"00",x"0f",x"ce"),
  1651 => (x"00",x"00",x"2a",x"16"),
  1652 => (x"00",x"00",x"00",x"00"),
  1653 => (x"00",x"00",x"0f",x"ce"),
  1654 => (x"00",x"00",x"2a",x"34"),
  1655 => (x"00",x"00",x"00",x"00"),
  1656 => (x"00",x"00",x"13",x"24"),
  1657 => (x"00",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"00",x"00",x"10",x"c8"),
  1660 => (x"00",x"00",x"00",x"00"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"00",x"00",x"10",x"94"),
  1663 => (x"db",x"86",x"fc",x"1e"),
  1664 => (x"fc",x"7e",x"70",x"87"),
  1665 => (x"1e",x"4f",x"26",x"8e"),
  1666 => (x"c0",x"48",x"f0",x"fe"),
  1667 => (x"79",x"09",x"cd",x"78"),
  1668 => (x"1e",x"4f",x"26",x"09"),
  1669 => (x"49",x"fc",x"e7",x"c1"),
  1670 => (x"4f",x"26",x"87",x"ed"),
  1671 => (x"bf",x"f0",x"fe",x"1e"),
  1672 => (x"1e",x"4f",x"26",x"48"),
  1673 => (x"c1",x"48",x"f0",x"fe"),
  1674 => (x"1e",x"4f",x"26",x"78"),
  1675 => (x"c0",x"48",x"f0",x"fe"),
  1676 => (x"1e",x"4f",x"26",x"78"),
  1677 => (x"52",x"c0",x"4a",x"71"),
  1678 => (x"0e",x"4f",x"26",x"51"),
  1679 => (x"5d",x"5c",x"5b",x"5e"),
  1680 => (x"71",x"86",x"f4",x"0e"),
  1681 => (x"7e",x"6d",x"97",x"4d"),
  1682 => (x"97",x"4c",x"a5",x"c1"),
  1683 => (x"a6",x"c8",x"48",x"6c"),
  1684 => (x"c4",x"48",x"6e",x"58"),
  1685 => (x"c5",x"05",x"a8",x"66"),
  1686 => (x"c0",x"48",x"ff",x"87"),
  1687 => (x"ca",x"ff",x"87",x"e6"),
  1688 => (x"49",x"a5",x"c2",x"87"),
  1689 => (x"71",x"4b",x"6c",x"97"),
  1690 => (x"6b",x"97",x"4b",x"a3"),
  1691 => (x"7e",x"6c",x"97",x"4b"),
  1692 => (x"80",x"c1",x"48",x"6e"),
  1693 => (x"c7",x"58",x"a6",x"c8"),
  1694 => (x"58",x"a6",x"cc",x"98"),
  1695 => (x"fe",x"7c",x"97",x"70"),
  1696 => (x"48",x"73",x"87",x"e1"),
  1697 => (x"4d",x"26",x"8e",x"f4"),
  1698 => (x"4b",x"26",x"4c",x"26"),
  1699 => (x"5e",x"0e",x"4f",x"26"),
  1700 => (x"f4",x"0e",x"5c",x"5b"),
  1701 => (x"d8",x"4c",x"71",x"86"),
  1702 => (x"ff",x"c3",x"4a",x"66"),
  1703 => (x"4b",x"a4",x"c2",x"9a"),
  1704 => (x"73",x"49",x"6c",x"97"),
  1705 => (x"51",x"72",x"49",x"a1"),
  1706 => (x"6e",x"7e",x"6c",x"97"),
  1707 => (x"c8",x"80",x"c1",x"48"),
  1708 => (x"98",x"c7",x"58",x"a6"),
  1709 => (x"70",x"58",x"a6",x"cc"),
  1710 => (x"26",x"8e",x"f4",x"54"),
  1711 => (x"26",x"4b",x"26",x"4c"),
  1712 => (x"86",x"fc",x"1e",x"4f"),
  1713 => (x"e0",x"87",x"e4",x"fd"),
  1714 => (x"c0",x"49",x"4a",x"bf"),
  1715 => (x"02",x"99",x"c0",x"e0"),
  1716 => (x"1e",x"72",x"87",x"cb"),
  1717 => (x"49",x"e8",x"e9",x"c2"),
  1718 => (x"c4",x"87",x"f3",x"fe"),
  1719 => (x"87",x"fc",x"fc",x"86"),
  1720 => (x"fe",x"fc",x"7e",x"70"),
  1721 => (x"26",x"8e",x"fc",x"87"),
  1722 => (x"e9",x"c2",x"1e",x"4f"),
  1723 => (x"c2",x"fd",x"49",x"e8"),
  1724 => (x"c1",x"eb",x"c1",x"87"),
  1725 => (x"87",x"cf",x"fc",x"49"),
  1726 => (x"26",x"87",x"ed",x"c4"),
  1727 => (x"5b",x"5e",x"0e",x"4f"),
  1728 => (x"fc",x"0e",x"5d",x"5c"),
  1729 => (x"ff",x"7e",x"71",x"86"),
  1730 => (x"e9",x"c2",x"4d",x"d4"),
  1731 => (x"ea",x"fc",x"49",x"e8"),
  1732 => (x"c0",x"4b",x"70",x"87"),
  1733 => (x"c2",x"04",x"ab",x"b7"),
  1734 => (x"f0",x"c3",x"87",x"f8"),
  1735 => (x"87",x"c9",x"05",x"ab"),
  1736 => (x"48",x"e0",x"ef",x"c1"),
  1737 => (x"d9",x"c2",x"78",x"c1"),
  1738 => (x"ab",x"e0",x"c3",x"87"),
  1739 => (x"c1",x"87",x"c9",x"05"),
  1740 => (x"c1",x"48",x"e4",x"ef"),
  1741 => (x"87",x"ca",x"c2",x"78"),
  1742 => (x"bf",x"e4",x"ef",x"c1"),
  1743 => (x"c2",x"87",x"c6",x"02"),
  1744 => (x"c2",x"4c",x"a3",x"c0"),
  1745 => (x"c1",x"4c",x"73",x"87"),
  1746 => (x"02",x"bf",x"e0",x"ef"),
  1747 => (x"74",x"87",x"e0",x"c0"),
  1748 => (x"29",x"b7",x"c4",x"49"),
  1749 => (x"e8",x"ef",x"c1",x"91"),
  1750 => (x"cf",x"4a",x"74",x"81"),
  1751 => (x"c1",x"92",x"c2",x"9a"),
  1752 => (x"70",x"30",x"72",x"48"),
  1753 => (x"72",x"ba",x"ff",x"4a"),
  1754 => (x"70",x"98",x"69",x"48"),
  1755 => (x"74",x"87",x"db",x"79"),
  1756 => (x"29",x"b7",x"c4",x"49"),
  1757 => (x"e8",x"ef",x"c1",x"91"),
  1758 => (x"cf",x"4a",x"74",x"81"),
  1759 => (x"c3",x"92",x"c2",x"9a"),
  1760 => (x"70",x"30",x"72",x"48"),
  1761 => (x"b0",x"69",x"48",x"4a"),
  1762 => (x"05",x"6e",x"79",x"70"),
  1763 => (x"ff",x"87",x"e7",x"c0"),
  1764 => (x"e1",x"c8",x"48",x"d0"),
  1765 => (x"c1",x"7d",x"c5",x"78"),
  1766 => (x"02",x"bf",x"e4",x"ef"),
  1767 => (x"e0",x"c3",x"87",x"c3"),
  1768 => (x"e0",x"ef",x"c1",x"7d"),
  1769 => (x"87",x"c3",x"02",x"bf"),
  1770 => (x"73",x"7d",x"f0",x"c3"),
  1771 => (x"48",x"d0",x"ff",x"7d"),
  1772 => (x"c0",x"78",x"e1",x"c8"),
  1773 => (x"ef",x"c1",x"78",x"e0"),
  1774 => (x"78",x"c0",x"48",x"e4"),
  1775 => (x"48",x"e0",x"ef",x"c1"),
  1776 => (x"e9",x"c2",x"78",x"c0"),
  1777 => (x"f2",x"f9",x"49",x"e8"),
  1778 => (x"c0",x"4b",x"70",x"87"),
  1779 => (x"fd",x"03",x"ab",x"b7"),
  1780 => (x"48",x"c0",x"87",x"c8"),
  1781 => (x"4d",x"26",x"8e",x"fc"),
  1782 => (x"4b",x"26",x"4c",x"26"),
  1783 => (x"00",x"00",x"4f",x"26"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"72",x"4a",x"c0",x"1e"),
  1803 => (x"c1",x"91",x"c4",x"49"),
  1804 => (x"c0",x"81",x"e8",x"ef"),
  1805 => (x"d0",x"82",x"c1",x"79"),
  1806 => (x"ee",x"04",x"aa",x"b7"),
  1807 => (x"0e",x"4f",x"26",x"87"),
  1808 => (x"5d",x"5c",x"5b",x"5e"),
  1809 => (x"f7",x"4d",x"71",x"0e"),
  1810 => (x"4a",x"75",x"87",x"e1"),
  1811 => (x"92",x"2a",x"b7",x"c4"),
  1812 => (x"82",x"e8",x"ef",x"c1"),
  1813 => (x"9c",x"cf",x"4c",x"75"),
  1814 => (x"49",x"6a",x"94",x"c2"),
  1815 => (x"c3",x"2b",x"74",x"4b"),
  1816 => (x"74",x"48",x"c2",x"9b"),
  1817 => (x"ff",x"4c",x"70",x"30"),
  1818 => (x"71",x"48",x"74",x"bc"),
  1819 => (x"f6",x"7a",x"70",x"98"),
  1820 => (x"48",x"73",x"87",x"f1"),
  1821 => (x"4c",x"26",x"4d",x"26"),
  1822 => (x"4f",x"26",x"4b",x"26"),
  1823 => (x"48",x"d0",x"ff",x"1e"),
  1824 => (x"71",x"78",x"e1",x"c8"),
  1825 => (x"08",x"d4",x"ff",x"48"),
  1826 => (x"48",x"66",x"c4",x"78"),
  1827 => (x"78",x"08",x"d4",x"ff"),
  1828 => (x"71",x"1e",x"4f",x"26"),
  1829 => (x"49",x"66",x"c4",x"4a"),
  1830 => (x"ff",x"49",x"72",x"1e"),
  1831 => (x"d0",x"ff",x"87",x"de"),
  1832 => (x"78",x"e0",x"c0",x"48"),
  1833 => (x"4f",x"26",x"8e",x"fc"),
  1834 => (x"71",x"1e",x"73",x"1e"),
  1835 => (x"49",x"66",x"c8",x"4b"),
  1836 => (x"c1",x"4a",x"73",x"1e"),
  1837 => (x"ff",x"49",x"a2",x"e0"),
  1838 => (x"8e",x"fc",x"87",x"d8"),
  1839 => (x"4f",x"26",x"4b",x"26"),
  1840 => (x"48",x"d0",x"ff",x"1e"),
  1841 => (x"71",x"78",x"c9",x"c8"),
  1842 => (x"08",x"d4",x"ff",x"48"),
  1843 => (x"1e",x"4f",x"26",x"78"),
  1844 => (x"eb",x"49",x"4a",x"71"),
  1845 => (x"48",x"d0",x"ff",x"87"),
  1846 => (x"4f",x"26",x"78",x"c8"),
  1847 => (x"71",x"1e",x"73",x"1e"),
  1848 => (x"c0",x"ea",x"c2",x"4b"),
  1849 => (x"87",x"c3",x"02",x"bf"),
  1850 => (x"ff",x"87",x"eb",x"c2"),
  1851 => (x"c9",x"c8",x"48",x"d0"),
  1852 => (x"c0",x"48",x"73",x"78"),
  1853 => (x"d4",x"ff",x"b0",x"e0"),
  1854 => (x"e9",x"c2",x"78",x"08"),
  1855 => (x"78",x"c0",x"48",x"f4"),
  1856 => (x"c5",x"02",x"66",x"c8"),
  1857 => (x"49",x"ff",x"c3",x"87"),
  1858 => (x"49",x"c0",x"87",x"c2"),
  1859 => (x"59",x"fc",x"e9",x"c2"),
  1860 => (x"c6",x"02",x"66",x"cc"),
  1861 => (x"d5",x"d5",x"c5",x"87"),
  1862 => (x"cf",x"87",x"c4",x"4a"),
  1863 => (x"c2",x"4a",x"ff",x"ff"),
  1864 => (x"c2",x"5a",x"c0",x"ea"),
  1865 => (x"c1",x"48",x"c0",x"ea"),
  1866 => (x"26",x"4b",x"26",x"78"),
  1867 => (x"5b",x"5e",x"0e",x"4f"),
  1868 => (x"71",x"0e",x"5d",x"5c"),
  1869 => (x"fc",x"e9",x"c2",x"4d"),
  1870 => (x"9d",x"75",x"4b",x"bf"),
  1871 => (x"49",x"87",x"cb",x"02"),
  1872 => (x"f3",x"c1",x"91",x"c8"),
  1873 => (x"82",x"71",x"4a",x"d4"),
  1874 => (x"f7",x"c1",x"87",x"c4"),
  1875 => (x"4c",x"c0",x"4a",x"d4"),
  1876 => (x"99",x"73",x"49",x"12"),
  1877 => (x"bf",x"f8",x"e9",x"c2"),
  1878 => (x"ff",x"b8",x"71",x"48"),
  1879 => (x"c1",x"78",x"08",x"d4"),
  1880 => (x"c8",x"84",x"2b",x"b7"),
  1881 => (x"e7",x"04",x"ac",x"b7"),
  1882 => (x"f4",x"e9",x"c2",x"87"),
  1883 => (x"80",x"c8",x"48",x"bf"),
  1884 => (x"58",x"f8",x"e9",x"c2"),
  1885 => (x"4c",x"26",x"4d",x"26"),
  1886 => (x"4f",x"26",x"4b",x"26"),
  1887 => (x"71",x"1e",x"73",x"1e"),
  1888 => (x"9a",x"4a",x"13",x"4b"),
  1889 => (x"72",x"87",x"cb",x"02"),
  1890 => (x"87",x"e1",x"fe",x"49"),
  1891 => (x"05",x"9a",x"4a",x"13"),
  1892 => (x"4b",x"26",x"87",x"f5"),
  1893 => (x"c2",x"1e",x"4f",x"26"),
  1894 => (x"49",x"bf",x"f4",x"e9"),
  1895 => (x"48",x"f4",x"e9",x"c2"),
  1896 => (x"c4",x"78",x"a1",x"c1"),
  1897 => (x"03",x"a9",x"b7",x"c0"),
  1898 => (x"d4",x"ff",x"87",x"db"),
  1899 => (x"f8",x"e9",x"c2",x"48"),
  1900 => (x"e9",x"c2",x"78",x"bf"),
  1901 => (x"c2",x"49",x"bf",x"f4"),
  1902 => (x"c1",x"48",x"f4",x"e9"),
  1903 => (x"c0",x"c4",x"78",x"a1"),
  1904 => (x"e5",x"04",x"a9",x"b7"),
  1905 => (x"48",x"d0",x"ff",x"87"),
  1906 => (x"ea",x"c2",x"78",x"c8"),
  1907 => (x"78",x"c0",x"48",x"c0"),
  1908 => (x"00",x"00",x"4f",x"26"),
  1909 => (x"00",x"00",x"00",x"00"),
  1910 => (x"00",x"00",x"00",x"00"),
  1911 => (x"5f",x"00",x"00",x"00"),
  1912 => (x"00",x"00",x"00",x"5f"),
  1913 => (x"00",x"03",x"03",x"00"),
  1914 => (x"00",x"00",x"03",x"03"),
  1915 => (x"14",x"7f",x"7f",x"14"),
  1916 => (x"00",x"14",x"7f",x"7f"),
  1917 => (x"6b",x"2e",x"24",x"00"),
  1918 => (x"00",x"12",x"3a",x"6b"),
  1919 => (x"18",x"36",x"6a",x"4c"),
  1920 => (x"00",x"32",x"56",x"6c"),
  1921 => (x"59",x"4f",x"7e",x"30"),
  1922 => (x"40",x"68",x"3a",x"77"),
  1923 => (x"07",x"04",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"03"),
  1925 => (x"3e",x"1c",x"00",x"00"),
  1926 => (x"00",x"00",x"41",x"63"),
  1927 => (x"63",x"41",x"00",x"00"),
  1928 => (x"00",x"00",x"1c",x"3e"),
  1929 => (x"1c",x"3e",x"2a",x"08"),
  1930 => (x"08",x"2a",x"3e",x"1c"),
  1931 => (x"3e",x"08",x"08",x"00"),
  1932 => (x"00",x"08",x"08",x"3e"),
  1933 => (x"e0",x"80",x"00",x"00"),
  1934 => (x"00",x"00",x"00",x"60"),
  1935 => (x"08",x"08",x"08",x"00"),
  1936 => (x"00",x"08",x"08",x"08"),
  1937 => (x"60",x"00",x"00",x"00"),
  1938 => (x"00",x"00",x"00",x"60"),
  1939 => (x"18",x"30",x"60",x"40"),
  1940 => (x"01",x"03",x"06",x"0c"),
  1941 => (x"59",x"7f",x"3e",x"00"),
  1942 => (x"00",x"3e",x"7f",x"4d"),
  1943 => (x"7f",x"06",x"04",x"00"),
  1944 => (x"00",x"00",x"00",x"7f"),
  1945 => (x"71",x"63",x"42",x"00"),
  1946 => (x"00",x"46",x"4f",x"59"),
  1947 => (x"49",x"63",x"22",x"00"),
  1948 => (x"00",x"36",x"7f",x"49"),
  1949 => (x"13",x"16",x"1c",x"18"),
  1950 => (x"00",x"10",x"7f",x"7f"),
  1951 => (x"45",x"67",x"27",x"00"),
  1952 => (x"00",x"39",x"7d",x"45"),
  1953 => (x"4b",x"7e",x"3c",x"00"),
  1954 => (x"00",x"30",x"79",x"49"),
  1955 => (x"71",x"01",x"01",x"00"),
  1956 => (x"00",x"07",x"0f",x"79"),
  1957 => (x"49",x"7f",x"36",x"00"),
  1958 => (x"00",x"36",x"7f",x"49"),
  1959 => (x"49",x"4f",x"06",x"00"),
  1960 => (x"00",x"1e",x"3f",x"69"),
  1961 => (x"66",x"00",x"00",x"00"),
  1962 => (x"00",x"00",x"00",x"66"),
  1963 => (x"e6",x"80",x"00",x"00"),
  1964 => (x"00",x"00",x"00",x"66"),
  1965 => (x"14",x"08",x"08",x"00"),
  1966 => (x"00",x"22",x"22",x"14"),
  1967 => (x"14",x"14",x"14",x"00"),
  1968 => (x"00",x"14",x"14",x"14"),
  1969 => (x"14",x"22",x"22",x"00"),
  1970 => (x"00",x"08",x"08",x"14"),
  1971 => (x"51",x"03",x"02",x"00"),
  1972 => (x"00",x"06",x"0f",x"59"),
  1973 => (x"5d",x"41",x"7f",x"3e"),
  1974 => (x"00",x"1e",x"1f",x"55"),
  1975 => (x"09",x"7f",x"7e",x"00"),
  1976 => (x"00",x"7e",x"7f",x"09"),
  1977 => (x"49",x"7f",x"7f",x"00"),
  1978 => (x"00",x"36",x"7f",x"49"),
  1979 => (x"63",x"3e",x"1c",x"00"),
  1980 => (x"00",x"41",x"41",x"41"),
  1981 => (x"41",x"7f",x"7f",x"00"),
  1982 => (x"00",x"1c",x"3e",x"63"),
  1983 => (x"49",x"7f",x"7f",x"00"),
  1984 => (x"00",x"41",x"41",x"49"),
  1985 => (x"09",x"7f",x"7f",x"00"),
  1986 => (x"00",x"01",x"01",x"09"),
  1987 => (x"41",x"7f",x"3e",x"00"),
  1988 => (x"00",x"7a",x"7b",x"49"),
  1989 => (x"08",x"7f",x"7f",x"00"),
  1990 => (x"00",x"7f",x"7f",x"08"),
  1991 => (x"7f",x"41",x"00",x"00"),
  1992 => (x"00",x"00",x"41",x"7f"),
  1993 => (x"40",x"60",x"20",x"00"),
  1994 => (x"00",x"3f",x"7f",x"40"),
  1995 => (x"1c",x"08",x"7f",x"7f"),
  1996 => (x"00",x"41",x"63",x"36"),
  1997 => (x"40",x"7f",x"7f",x"00"),
  1998 => (x"00",x"40",x"40",x"40"),
  1999 => (x"0c",x"06",x"7f",x"7f"),
  2000 => (x"00",x"7f",x"7f",x"06"),
  2001 => (x"0c",x"06",x"7f",x"7f"),
  2002 => (x"00",x"7f",x"7f",x"18"),
  2003 => (x"41",x"7f",x"3e",x"00"),
  2004 => (x"00",x"3e",x"7f",x"41"),
  2005 => (x"09",x"7f",x"7f",x"00"),
  2006 => (x"00",x"06",x"0f",x"09"),
  2007 => (x"61",x"41",x"7f",x"3e"),
  2008 => (x"00",x"40",x"7e",x"7f"),
  2009 => (x"09",x"7f",x"7f",x"00"),
  2010 => (x"00",x"66",x"7f",x"19"),
  2011 => (x"4d",x"6f",x"26",x"00"),
  2012 => (x"00",x"32",x"7b",x"59"),
  2013 => (x"7f",x"01",x"01",x"00"),
  2014 => (x"00",x"01",x"01",x"7f"),
  2015 => (x"40",x"7f",x"3f",x"00"),
  2016 => (x"00",x"3f",x"7f",x"40"),
  2017 => (x"70",x"3f",x"0f",x"00"),
  2018 => (x"00",x"0f",x"3f",x"70"),
  2019 => (x"18",x"30",x"7f",x"7f"),
  2020 => (x"00",x"7f",x"7f",x"30"),
  2021 => (x"1c",x"36",x"63",x"41"),
  2022 => (x"41",x"63",x"36",x"1c"),
  2023 => (x"7c",x"06",x"03",x"01"),
  2024 => (x"01",x"03",x"06",x"7c"),
  2025 => (x"4d",x"59",x"71",x"61"),
  2026 => (x"00",x"41",x"43",x"47"),
  2027 => (x"7f",x"7f",x"00",x"00"),
  2028 => (x"00",x"00",x"41",x"41"),
  2029 => (x"0c",x"06",x"03",x"01"),
  2030 => (x"40",x"60",x"30",x"18"),
  2031 => (x"41",x"41",x"00",x"00"),
  2032 => (x"00",x"00",x"7f",x"7f"),
  2033 => (x"03",x"06",x"0c",x"08"),
  2034 => (x"00",x"08",x"0c",x"06"),
  2035 => (x"80",x"80",x"80",x"80"),
  2036 => (x"00",x"80",x"80",x"80"),
  2037 => (x"03",x"00",x"00",x"00"),
  2038 => (x"00",x"00",x"04",x"07"),
  2039 => (x"54",x"74",x"20",x"00"),
  2040 => (x"00",x"78",x"7c",x"54"),
  2041 => (x"44",x"7f",x"7f",x"00"),
  2042 => (x"00",x"38",x"7c",x"44"),
  2043 => (x"44",x"7c",x"38",x"00"),
  2044 => (x"00",x"00",x"44",x"44"),
  2045 => (x"44",x"7c",x"38",x"00"),
  2046 => (x"00",x"7f",x"7f",x"44"),
  2047 => (x"54",x"7c",x"38",x"00"),
  2048 => (x"00",x"18",x"5c",x"54"),
  2049 => (x"7f",x"7e",x"04",x"00"),
  2050 => (x"00",x"00",x"05",x"05"),
  2051 => (x"a4",x"bc",x"18",x"00"),
  2052 => (x"00",x"7c",x"fc",x"a4"),
  2053 => (x"04",x"7f",x"7f",x"00"),
  2054 => (x"00",x"78",x"7c",x"04"),
  2055 => (x"3d",x"00",x"00",x"00"),
  2056 => (x"00",x"00",x"40",x"7d"),
  2057 => (x"80",x"80",x"80",x"00"),
  2058 => (x"00",x"00",x"7d",x"fd"),
  2059 => (x"10",x"7f",x"7f",x"00"),
  2060 => (x"00",x"44",x"6c",x"38"),
  2061 => (x"3f",x"00",x"00",x"00"),
  2062 => (x"00",x"00",x"40",x"7f"),
  2063 => (x"18",x"0c",x"7c",x"7c"),
  2064 => (x"00",x"78",x"7c",x"0c"),
  2065 => (x"04",x"7c",x"7c",x"00"),
  2066 => (x"00",x"78",x"7c",x"04"),
  2067 => (x"44",x"7c",x"38",x"00"),
  2068 => (x"00",x"38",x"7c",x"44"),
  2069 => (x"24",x"fc",x"fc",x"00"),
  2070 => (x"00",x"18",x"3c",x"24"),
  2071 => (x"24",x"3c",x"18",x"00"),
  2072 => (x"00",x"fc",x"fc",x"24"),
  2073 => (x"04",x"7c",x"7c",x"00"),
  2074 => (x"00",x"08",x"0c",x"04"),
  2075 => (x"54",x"5c",x"48",x"00"),
  2076 => (x"00",x"20",x"74",x"54"),
  2077 => (x"7f",x"3f",x"04",x"00"),
  2078 => (x"00",x"00",x"44",x"44"),
  2079 => (x"40",x"7c",x"3c",x"00"),
  2080 => (x"00",x"7c",x"7c",x"40"),
  2081 => (x"60",x"3c",x"1c",x"00"),
  2082 => (x"00",x"1c",x"3c",x"60"),
  2083 => (x"30",x"60",x"7c",x"3c"),
  2084 => (x"00",x"3c",x"7c",x"60"),
  2085 => (x"10",x"38",x"6c",x"44"),
  2086 => (x"00",x"44",x"6c",x"38"),
  2087 => (x"e0",x"bc",x"1c",x"00"),
  2088 => (x"00",x"1c",x"3c",x"60"),
  2089 => (x"74",x"64",x"44",x"00"),
  2090 => (x"00",x"44",x"4c",x"5c"),
  2091 => (x"3e",x"08",x"08",x"00"),
  2092 => (x"00",x"41",x"41",x"77"),
  2093 => (x"7f",x"00",x"00",x"00"),
  2094 => (x"00",x"00",x"00",x"7f"),
  2095 => (x"77",x"41",x"41",x"00"),
  2096 => (x"00",x"08",x"08",x"3e"),
  2097 => (x"03",x"01",x"01",x"02"),
  2098 => (x"00",x"01",x"02",x"02"),
  2099 => (x"7f",x"7f",x"7f",x"7f"),
  2100 => (x"00",x"7f",x"7f",x"7f"),
  2101 => (x"1c",x"1c",x"08",x"08"),
  2102 => (x"7f",x"7f",x"3e",x"3e"),
  2103 => (x"3e",x"3e",x"7f",x"7f"),
  2104 => (x"08",x"08",x"1c",x"1c"),
  2105 => (x"7c",x"18",x"10",x"00"),
  2106 => (x"00",x"10",x"18",x"7c"),
  2107 => (x"7c",x"30",x"10",x"00"),
  2108 => (x"00",x"10",x"30",x"7c"),
  2109 => (x"60",x"60",x"30",x"10"),
  2110 => (x"00",x"06",x"1e",x"78"),
  2111 => (x"18",x"3c",x"66",x"42"),
  2112 => (x"00",x"42",x"66",x"3c"),
  2113 => (x"c2",x"6a",x"38",x"78"),
  2114 => (x"00",x"38",x"6c",x"c6"),
  2115 => (x"60",x"00",x"00",x"60"),
  2116 => (x"00",x"60",x"00",x"00"),
  2117 => (x"5c",x"5b",x"5e",x"0e"),
  2118 => (x"86",x"fc",x"0e",x"5d"),
  2119 => (x"ea",x"c2",x"7e",x"71"),
  2120 => (x"c0",x"4c",x"bf",x"c8"),
  2121 => (x"c4",x"1e",x"c0",x"4b"),
  2122 => (x"c4",x"02",x"ab",x"66"),
  2123 => (x"c2",x"4d",x"c0",x"87"),
  2124 => (x"75",x"4d",x"c1",x"87"),
  2125 => (x"ee",x"49",x"73",x"1e"),
  2126 => (x"86",x"c8",x"87",x"e2"),
  2127 => (x"ef",x"49",x"e0",x"c0"),
  2128 => (x"a4",x"c4",x"87",x"eb"),
  2129 => (x"f0",x"49",x"6a",x"4a"),
  2130 => (x"c9",x"f1",x"87",x"f2"),
  2131 => (x"c1",x"84",x"cc",x"87"),
  2132 => (x"ab",x"b7",x"c8",x"83"),
  2133 => (x"87",x"cd",x"ff",x"04"),
  2134 => (x"4d",x"26",x"8e",x"fc"),
  2135 => (x"4b",x"26",x"4c",x"26"),
  2136 => (x"71",x"1e",x"4f",x"26"),
  2137 => (x"cc",x"ea",x"c2",x"4a"),
  2138 => (x"cc",x"ea",x"c2",x"5a"),
  2139 => (x"49",x"78",x"c7",x"48"),
  2140 => (x"26",x"87",x"e1",x"fe"),
  2141 => (x"1e",x"73",x"1e",x"4f"),
  2142 => (x"b7",x"c0",x"4a",x"71"),
  2143 => (x"87",x"d3",x"03",x"aa"),
  2144 => (x"bf",x"f0",x"d4",x"c2"),
  2145 => (x"c1",x"87",x"c4",x"05"),
  2146 => (x"c0",x"87",x"c2",x"4b"),
  2147 => (x"f4",x"d4",x"c2",x"4b"),
  2148 => (x"c2",x"87",x"c4",x"5b"),
  2149 => (x"fc",x"5a",x"f4",x"d4"),
  2150 => (x"f0",x"d4",x"c2",x"48"),
  2151 => (x"c1",x"4a",x"78",x"bf"),
  2152 => (x"a2",x"c0",x"c1",x"9a"),
  2153 => (x"87",x"e7",x"ec",x"49"),
  2154 => (x"4f",x"26",x"4b",x"26"),
  2155 => (x"c4",x"4a",x"71",x"1e"),
  2156 => (x"49",x"72",x"1e",x"66"),
  2157 => (x"fc",x"87",x"f1",x"eb"),
  2158 => (x"1e",x"4f",x"26",x"8e"),
  2159 => (x"c3",x"48",x"d4",x"ff"),
  2160 => (x"d0",x"ff",x"78",x"ff"),
  2161 => (x"78",x"e1",x"c0",x"48"),
  2162 => (x"c1",x"48",x"d4",x"ff"),
  2163 => (x"c4",x"48",x"71",x"78"),
  2164 => (x"08",x"d4",x"ff",x"30"),
  2165 => (x"48",x"d0",x"ff",x"78"),
  2166 => (x"26",x"78",x"e0",x"c0"),
  2167 => (x"5b",x"5e",x"0e",x"4f"),
  2168 => (x"f0",x"0e",x"5d",x"5c"),
  2169 => (x"48",x"a6",x"c8",x"86"),
  2170 => (x"bf",x"ec",x"78",x"c0"),
  2171 => (x"c2",x"80",x"fc",x"7e"),
  2172 => (x"78",x"bf",x"c8",x"ea"),
  2173 => (x"bf",x"d0",x"ea",x"c2"),
  2174 => (x"4c",x"bf",x"e8",x"4d"),
  2175 => (x"bf",x"f0",x"d4",x"c2"),
  2176 => (x"87",x"f9",x"e3",x"49"),
  2177 => (x"f6",x"e8",x"49",x"c7"),
  2178 => (x"c2",x"49",x"70",x"87"),
  2179 => (x"87",x"cf",x"05",x"99"),
  2180 => (x"bf",x"e8",x"d4",x"c2"),
  2181 => (x"6e",x"b9",x"ff",x"49"),
  2182 => (x"02",x"99",x"c1",x"99"),
  2183 => (x"cb",x"87",x"c0",x"c2"),
  2184 => (x"cf",x"cc",x"49",x"ee"),
  2185 => (x"58",x"a6",x"d0",x"87"),
  2186 => (x"d2",x"e8",x"49",x"c7"),
  2187 => (x"05",x"98",x"70",x"87"),
  2188 => (x"49",x"6e",x"87",x"c8"),
  2189 => (x"c1",x"02",x"99",x"c1"),
  2190 => (x"66",x"cc",x"87",x"c2"),
  2191 => (x"7e",x"bf",x"ec",x"4b"),
  2192 => (x"bf",x"f0",x"d4",x"c2"),
  2193 => (x"87",x"f5",x"e2",x"49"),
  2194 => (x"f3",x"cb",x"49",x"73"),
  2195 => (x"02",x"98",x"70",x"87"),
  2196 => (x"d4",x"c2",x"87",x"d7"),
  2197 => (x"c1",x"49",x"bf",x"d0"),
  2198 => (x"d4",x"d4",x"c2",x"b9"),
  2199 => (x"da",x"fd",x"71",x"59"),
  2200 => (x"49",x"ee",x"cb",x"87"),
  2201 => (x"70",x"87",x"cd",x"cb"),
  2202 => (x"e7",x"49",x"c7",x"4b"),
  2203 => (x"98",x"70",x"87",x"d1"),
  2204 => (x"87",x"c9",x"ff",x"05"),
  2205 => (x"99",x"c1",x"49",x"6e"),
  2206 => (x"87",x"c1",x"ff",x"05"),
  2207 => (x"bf",x"f0",x"d4",x"c2"),
  2208 => (x"c2",x"ba",x"c1",x"4a"),
  2209 => (x"fc",x"5a",x"f4",x"d4"),
  2210 => (x"c1",x"0a",x"7a",x"0a"),
  2211 => (x"a2",x"c0",x"c1",x"9a"),
  2212 => (x"87",x"fb",x"e8",x"49"),
  2213 => (x"e6",x"49",x"da",x"c1"),
  2214 => (x"a6",x"c8",x"87",x"e5"),
  2215 => (x"c2",x"78",x"c1",x"48"),
  2216 => (x"6e",x"48",x"e8",x"d4"),
  2217 => (x"f0",x"d4",x"c2",x"78"),
  2218 => (x"c7",x"c1",x"05",x"bf"),
  2219 => (x"c0",x"c0",x"c8",x"87"),
  2220 => (x"c8",x"d7",x"c2",x"4b"),
  2221 => (x"49",x"15",x"4d",x"7e"),
  2222 => (x"87",x"c3",x"e6",x"49"),
  2223 => (x"c0",x"02",x"98",x"70"),
  2224 => (x"b4",x"73",x"87",x"c2"),
  2225 => (x"05",x"2b",x"b7",x"c1"),
  2226 => (x"74",x"87",x"eb",x"ff"),
  2227 => (x"99",x"ff",x"c3",x"49"),
  2228 => (x"49",x"c0",x"1e",x"71"),
  2229 => (x"74",x"87",x"d5",x"fb"),
  2230 => (x"29",x"b7",x"c8",x"49"),
  2231 => (x"49",x"c1",x"1e",x"71"),
  2232 => (x"c8",x"87",x"c9",x"fb"),
  2233 => (x"49",x"fd",x"c3",x"86"),
  2234 => (x"c3",x"87",x"d4",x"e5"),
  2235 => (x"ce",x"e5",x"49",x"fa"),
  2236 => (x"87",x"d1",x"c8",x"87"),
  2237 => (x"ff",x"c3",x"49",x"74"),
  2238 => (x"2c",x"b7",x"c8",x"99"),
  2239 => (x"9c",x"74",x"b4",x"71"),
  2240 => (x"ff",x"87",x"df",x"02"),
  2241 => (x"49",x"7e",x"bf",x"c8"),
  2242 => (x"bf",x"ec",x"d4",x"c2"),
  2243 => (x"a9",x"e0",x"c2",x"89"),
  2244 => (x"87",x"c5",x"c0",x"03"),
  2245 => (x"cf",x"c0",x"4c",x"c0"),
  2246 => (x"ec",x"d4",x"c2",x"87"),
  2247 => (x"c0",x"78",x"6e",x"48"),
  2248 => (x"d4",x"c2",x"87",x"c6"),
  2249 => (x"78",x"c0",x"48",x"ec"),
  2250 => (x"99",x"c8",x"49",x"74"),
  2251 => (x"87",x"ce",x"c0",x"05"),
  2252 => (x"e4",x"49",x"f5",x"c3"),
  2253 => (x"49",x"70",x"87",x"c9"),
  2254 => (x"c0",x"02",x"99",x"c2"),
  2255 => (x"ea",x"c2",x"87",x"ea"),
  2256 => (x"c0",x"02",x"bf",x"cc"),
  2257 => (x"c1",x"48",x"87",x"ca"),
  2258 => (x"d0",x"ea",x"c2",x"88"),
  2259 => (x"87",x"d3",x"c0",x"58"),
  2260 => (x"c1",x"48",x"66",x"c4"),
  2261 => (x"7e",x"70",x"80",x"e0"),
  2262 => (x"c0",x"02",x"bf",x"6e"),
  2263 => (x"ff",x"4b",x"87",x"c5"),
  2264 => (x"c8",x"0f",x"73",x"49"),
  2265 => (x"78",x"c1",x"48",x"a6"),
  2266 => (x"99",x"c4",x"49",x"74"),
  2267 => (x"87",x"ce",x"c0",x"05"),
  2268 => (x"e3",x"49",x"f2",x"c3"),
  2269 => (x"49",x"70",x"87",x"c9"),
  2270 => (x"c0",x"02",x"99",x"c2"),
  2271 => (x"ea",x"c2",x"87",x"f0"),
  2272 => (x"48",x"7e",x"bf",x"cc"),
  2273 => (x"03",x"a8",x"b7",x"c7"),
  2274 => (x"6e",x"87",x"cb",x"c0"),
  2275 => (x"c2",x"80",x"c1",x"48"),
  2276 => (x"c0",x"58",x"d0",x"ea"),
  2277 => (x"66",x"c4",x"87",x"d3"),
  2278 => (x"80",x"e0",x"c1",x"48"),
  2279 => (x"bf",x"6e",x"7e",x"70"),
  2280 => (x"87",x"c5",x"c0",x"02"),
  2281 => (x"73",x"49",x"fe",x"4b"),
  2282 => (x"48",x"a6",x"c8",x"0f"),
  2283 => (x"fd",x"c3",x"78",x"c1"),
  2284 => (x"87",x"cb",x"e2",x"49"),
  2285 => (x"99",x"c2",x"49",x"70"),
  2286 => (x"87",x"e6",x"c0",x"02"),
  2287 => (x"bf",x"cc",x"ea",x"c2"),
  2288 => (x"87",x"c9",x"c0",x"02"),
  2289 => (x"48",x"cc",x"ea",x"c2"),
  2290 => (x"d0",x"c0",x"78",x"c0"),
  2291 => (x"4a",x"66",x"c4",x"87"),
  2292 => (x"6a",x"82",x"e0",x"c1"),
  2293 => (x"87",x"c5",x"c0",x"02"),
  2294 => (x"73",x"49",x"fd",x"4b"),
  2295 => (x"48",x"a6",x"c8",x"0f"),
  2296 => (x"fa",x"c3",x"78",x"c1"),
  2297 => (x"87",x"d7",x"e1",x"49"),
  2298 => (x"99",x"c2",x"49",x"70"),
  2299 => (x"87",x"ed",x"c0",x"02"),
  2300 => (x"bf",x"cc",x"ea",x"c2"),
  2301 => (x"a8",x"b7",x"c7",x"48"),
  2302 => (x"87",x"c9",x"c0",x"03"),
  2303 => (x"48",x"cc",x"ea",x"c2"),
  2304 => (x"d3",x"c0",x"78",x"c7"),
  2305 => (x"48",x"66",x"c4",x"87"),
  2306 => (x"70",x"80",x"e0",x"c1"),
  2307 => (x"02",x"bf",x"6e",x"7e"),
  2308 => (x"4b",x"87",x"c5",x"c0"),
  2309 => (x"0f",x"73",x"49",x"fc"),
  2310 => (x"c1",x"48",x"a6",x"c8"),
  2311 => (x"c3",x"48",x"74",x"78"),
  2312 => (x"7e",x"70",x"98",x"f0"),
  2313 => (x"c0",x"05",x"98",x"48"),
  2314 => (x"da",x"c1",x"87",x"ce"),
  2315 => (x"87",x"cf",x"e0",x"49"),
  2316 => (x"99",x"c2",x"49",x"70"),
  2317 => (x"87",x"d0",x"c2",x"02"),
  2318 => (x"c3",x"49",x"ee",x"cb"),
  2319 => (x"a6",x"d0",x"87",x"f6"),
  2320 => (x"c4",x"ea",x"c2",x"58"),
  2321 => (x"c2",x"50",x"c0",x"48"),
  2322 => (x"bf",x"97",x"c4",x"ea"),
  2323 => (x"87",x"d8",x"c1",x"05"),
  2324 => (x"cd",x"c0",x"05",x"6e"),
  2325 => (x"49",x"da",x"c1",x"87"),
  2326 => (x"87",x"e3",x"df",x"ff"),
  2327 => (x"c1",x"02",x"98",x"70"),
  2328 => (x"bf",x"e8",x"87",x"c6"),
  2329 => (x"ff",x"c3",x"49",x"4b"),
  2330 => (x"2b",x"b7",x"c8",x"99"),
  2331 => (x"d4",x"c2",x"b3",x"71"),
  2332 => (x"ff",x"49",x"bf",x"f0"),
  2333 => (x"cc",x"87",x"c6",x"da"),
  2334 => (x"c3",x"c3",x"49",x"66"),
  2335 => (x"02",x"98",x"70",x"87"),
  2336 => (x"c2",x"87",x"c6",x"c0"),
  2337 => (x"c1",x"48",x"c4",x"ea"),
  2338 => (x"c4",x"ea",x"c2",x"50"),
  2339 => (x"c0",x"05",x"bf",x"97"),
  2340 => (x"49",x"73",x"87",x"d6"),
  2341 => (x"05",x"99",x"f0",x"c3"),
  2342 => (x"c1",x"87",x"c7",x"ff"),
  2343 => (x"de",x"ff",x"49",x"da"),
  2344 => (x"98",x"70",x"87",x"dd"),
  2345 => (x"87",x"fa",x"fe",x"05"),
  2346 => (x"c2",x"48",x"a6",x"cc"),
  2347 => (x"78",x"bf",x"cc",x"ea"),
  2348 => (x"cc",x"49",x"66",x"cc"),
  2349 => (x"48",x"66",x"c4",x"91"),
  2350 => (x"7e",x"70",x"80",x"71"),
  2351 => (x"c0",x"02",x"bf",x"6e"),
  2352 => (x"cc",x"4b",x"87",x"c6"),
  2353 => (x"0f",x"73",x"49",x"66"),
  2354 => (x"c0",x"02",x"9d",x"75"),
  2355 => (x"02",x"6d",x"87",x"e9"),
  2356 => (x"6d",x"87",x"e4",x"c0"),
  2357 => (x"e6",x"dd",x"ff",x"49"),
  2358 => (x"c1",x"49",x"70",x"87"),
  2359 => (x"cb",x"c0",x"02",x"99"),
  2360 => (x"4b",x"a5",x"c4",x"87"),
  2361 => (x"bf",x"cc",x"ea",x"c2"),
  2362 => (x"0f",x"4b",x"6b",x"49"),
  2363 => (x"c0",x"02",x"85",x"c8"),
  2364 => (x"05",x"6d",x"87",x"c5"),
  2365 => (x"c8",x"87",x"dc",x"ff"),
  2366 => (x"c8",x"c0",x"02",x"66"),
  2367 => (x"cc",x"ea",x"c2",x"87"),
  2368 => (x"cf",x"f0",x"49",x"bf"),
  2369 => (x"26",x"8e",x"f0",x"87"),
  2370 => (x"26",x"4c",x"26",x"4d"),
  2371 => (x"00",x"4f",x"26",x"4b"),
  2372 => (x"00",x"00",x"00",x"00"),
  2373 => (x"00",x"00",x"00",x"10"),
  2374 => (x"14",x"11",x"12",x"58"),
  2375 => (x"23",x"1c",x"1b",x"1d"),
  2376 => (x"94",x"91",x"59",x"5a"),
  2377 => (x"f4",x"eb",x"f2",x"f5"),
  2378 => (x"00",x"00",x"00",x"00"),
  2379 => (x"00",x"00",x"00",x"00"),
  2380 => (x"00",x"00",x"00",x"00"),
  2381 => (x"ff",x"4a",x"71",x"1e"),
  2382 => (x"72",x"49",x"bf",x"c8"),
  2383 => (x"4f",x"26",x"48",x"a1"),
  2384 => (x"bf",x"c8",x"ff",x"1e"),
  2385 => (x"c0",x"c0",x"fe",x"89"),
  2386 => (x"a9",x"c0",x"c0",x"c0"),
  2387 => (x"c0",x"87",x"c4",x"01"),
  2388 => (x"c1",x"87",x"c2",x"4a"),
  2389 => (x"26",x"48",x"72",x"4a"),
  2390 => (x"1e",x"73",x"1e",x"4f"),
  2391 => (x"e6",x"c1",x"4b",x"c0"),
  2392 => (x"50",x"c0",x"48",x"c0"),
  2393 => (x"bf",x"d8",x"d7",x"c2"),
  2394 => (x"c1",x"e3",x"fe",x"49"),
  2395 => (x"05",x"98",x"70",x"87"),
  2396 => (x"d6",x"c2",x"87",x"c4"),
  2397 => (x"e6",x"c1",x"4b",x"cc"),
  2398 => (x"50",x"c1",x"48",x"c0"),
  2399 => (x"bf",x"dc",x"d7",x"c2"),
  2400 => (x"e9",x"e2",x"fe",x"49"),
  2401 => (x"26",x"48",x"73",x"87"),
  2402 => (x"00",x"4f",x"26",x"4b"),
  2403 => (x"5f",x"43",x"42",x"47"),
  2404 => (x"53",x"4f",x"49",x"42"),
  2405 => (x"4e",x"49",x"42",x"2e"),
  2406 => (x"74",x"6f",x"6e",x"20"),
  2407 => (x"75",x"6f",x"66",x"20"),
  2408 => (x"6f",x"20",x"64",x"6e"),
  2409 => (x"44",x"53",x"20",x"6e"),
  2410 => (x"72",x"61",x"63",x"20"),
  2411 => (x"00",x"00",x"00",x"64"),
  2412 => (x"5f",x"43",x"42",x"47"),
  2413 => (x"53",x"4f",x"49",x"42"),
  2414 => (x"00",x"4e",x"49",x"42"),
  2415 => (x"4f",x"54",x"55",x"41"),
  2416 => (x"54",x"4f",x"4f",x"42"),
  2417 => (x"00",x"00",x"42",x"47"),
  2418 => (x"11",x"14",x"12",x"58"),
  2419 => (x"23",x"1c",x"1b",x"1d"),
  2420 => (x"91",x"94",x"59",x"5a"),
  2421 => (x"f4",x"eb",x"f2",x"f5"),
  2422 => (x"00",x"00",x"25",x"b0"),
  2423 => (x"00",x"00",x"25",x"bc"),
  2424 => (x"00",x"00",x"1a",x"13"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

