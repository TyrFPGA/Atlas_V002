
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"fa",x"c2",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"dc",x"fa",x"c2"),
    14 => (x"48",x"e8",x"e7",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ea",x"e3"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"e8",x"e7"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"e7",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"e8"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"ec",x"e7",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"f0",x"e7",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"f0",x"e7",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"f0",x"e7"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"f7",x"e7"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"f8",x"e7"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"f9",x"e7",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"e7",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"f9"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"fa",x"e7",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"f5",x"e7"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"f6",x"e7",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"e7",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"f7"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"f8",x"e7",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"f0",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"d6"),
   330 => (x"1e",x"ce",x"e8",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"dd",x"f2",x"c0",x"7e"),
   337 => (x"e9",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"c4"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"d9",x"f2"),
   343 => (x"4a",x"e0",x"e9",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"ef",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"d4"),
   350 => (x"bf",x"9f",x"cc",x"f0"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"d4",x"ef",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"e8",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"ce"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"d9",x"f2"),
   365 => (x"4a",x"e0",x"e9",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"d6",x"f0"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"dd",x"f2"),
   372 => (x"4a",x"c4",x"e9",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"cc",x"f0",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"f0",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"cd"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"ce",x"e8",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"d9",x"e8",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"da",x"e8"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"db",x"e8",x"c2"),
   400 => (x"f0",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"d2"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"d6",x"f0"),
   404 => (x"bf",x"97",x"dc",x"e8"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"dd",x"e8"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"f4",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"e3"),
   410 => (x"97",x"de",x"e8",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"d6",x"f0",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"d9",x"f2",x"c0",x"87"),
   415 => (x"e9",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"e0"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"ce",x"f0"),
   422 => (x"5c",x"f7",x"f4",x"c2"),
   423 => (x"97",x"f3",x"e8",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"f2",x"e8",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"f4",x"e8",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"f5",x"e8"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"e3",x"f4",x"c2",x"91"),
   434 => (x"f4",x"c2",x"81",x"bf"),
   435 => (x"e8",x"c2",x"59",x"eb"),
   436 => (x"4a",x"bf",x"97",x"fb"),
   437 => (x"e8",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"fa"),
   439 => (x"e8",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"fc"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"fd",x"e8",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"f4",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"ef"),
   447 => (x"f4",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"ef"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"e0",x"e8",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"df",x"e8",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"f7",x"f4"),
   457 => (x"bf",x"97",x"e5",x"e8"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"e4",x"e8"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"f3",x"f4",x"c2"),
   463 => (x"48",x"eb",x"f4",x"c2"),
   464 => (x"f4",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"e7"),
   466 => (x"f7",x"f4",x"c2",x"78"),
   467 => (x"eb",x"f4",x"c2",x"48"),
   468 => (x"f4",x"c2",x"78",x"bf"),
   469 => (x"f4",x"c2",x"48",x"fb"),
   470 => (x"c2",x"78",x"bf",x"ef"),
   471 => (x"02",x"bf",x"d6",x"f0"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"f3",x"f4",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"da",x"f0",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"d6",x"f0"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"f4",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"e3"),
   492 => (x"ab",x"bf",x"d5",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"d9",x"f2"),
   495 => (x"73",x"1e",x"ce",x"e8"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"d6",x"f0",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"ce",x"e8"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"ce",x"e8",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c0",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"e9",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d3",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"de",x"f0",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d1",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"ce",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"d6",x"f0"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"48",x"6e",x"7e",x"c0"),
   556 => (x"80",x"bf",x"66",x"c4"),
   557 => (x"78",x"08",x"66",x"c4"),
   558 => (x"a4",x"cc",x"7c",x"c0"),
   559 => (x"bf",x"66",x"c4",x"49"),
   560 => (x"49",x"a4",x"d0",x"79"),
   561 => (x"48",x"c1",x"79",x"c0"),
   562 => (x"48",x"c0",x"87",x"c2"),
   563 => (x"ee",x"fa",x"8e",x"f8"),
   564 => (x"5b",x"5e",x"0e",x"87"),
   565 => (x"4c",x"71",x"0e",x"5c"),
   566 => (x"cb",x"c1",x"02",x"9c"),
   567 => (x"49",x"a4",x"c8",x"87"),
   568 => (x"c3",x"c1",x"02",x"69"),
   569 => (x"cc",x"49",x"6c",x"87"),
   570 => (x"80",x"71",x"48",x"66"),
   571 => (x"70",x"58",x"a6",x"d0"),
   572 => (x"d2",x"f0",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e5",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"ff",x"f9",x"49"),
   578 => (x"f0",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"ce"),
   580 => (x"cc",x"7c",x"71",x"81"),
   581 => (x"f0",x"c2",x"b9",x"66"),
   582 => (x"ff",x"4a",x"bf",x"d2"),
   583 => (x"71",x"99",x"72",x"ba"),
   584 => (x"db",x"ff",x"05",x"99"),
   585 => (x"7c",x"66",x"cc",x"87"),
   586 => (x"1e",x"87",x"d6",x"f9"),
   587 => (x"4b",x"71",x"1e",x"73"),
   588 => (x"87",x"c7",x"02",x"9b"),
   589 => (x"69",x"49",x"a3",x"c8"),
   590 => (x"c0",x"87",x"c5",x"05"),
   591 => (x"87",x"f6",x"c0",x"48"),
   592 => (x"bf",x"e7",x"f4",x"c2"),
   593 => (x"4a",x"a3",x"c4",x"49"),
   594 => (x"8a",x"c2",x"4a",x"6a"),
   595 => (x"bf",x"ce",x"f0",x"c2"),
   596 => (x"49",x"a1",x"72",x"92"),
   597 => (x"bf",x"d2",x"f0",x"c2"),
   598 => (x"72",x"9a",x"6b",x"4a"),
   599 => (x"f2",x"c0",x"49",x"a1"),
   600 => (x"66",x"c8",x"59",x"d9"),
   601 => (x"e6",x"ea",x"71",x"1e"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"87",x"c4",x"05",x"98"),
   604 => (x"87",x"c2",x"48",x"c0"),
   605 => (x"ca",x"f8",x"48",x"c1"),
   606 => (x"1e",x"73",x"1e",x"87"),
   607 => (x"02",x"9b",x"4b",x"71"),
   608 => (x"a3",x"c8",x"87",x"c7"),
   609 => (x"c5",x"05",x"69",x"49"),
   610 => (x"c0",x"48",x"c0",x"87"),
   611 => (x"f4",x"c2",x"87",x"f6"),
   612 => (x"c4",x"49",x"bf",x"e7"),
   613 => (x"4a",x"6a",x"4a",x"a3"),
   614 => (x"f0",x"c2",x"8a",x"c2"),
   615 => (x"72",x"92",x"bf",x"ce"),
   616 => (x"f0",x"c2",x"49",x"a1"),
   617 => (x"6b",x"4a",x"bf",x"d2"),
   618 => (x"49",x"a1",x"72",x"9a"),
   619 => (x"59",x"d9",x"f2",x"c0"),
   620 => (x"71",x"1e",x"66",x"c8"),
   621 => (x"c4",x"87",x"d1",x"e6"),
   622 => (x"05",x"98",x"70",x"86"),
   623 => (x"48",x"c0",x"87",x"c4"),
   624 => (x"48",x"c1",x"87",x"c2"),
   625 => (x"0e",x"87",x"fc",x"f6"),
   626 => (x"5d",x"5c",x"5b",x"5e"),
   627 => (x"4b",x"71",x"1e",x"0e"),
   628 => (x"73",x"4d",x"66",x"d4"),
   629 => (x"cc",x"c1",x"02",x"9b"),
   630 => (x"49",x"a3",x"c8",x"87"),
   631 => (x"c4",x"c1",x"02",x"69"),
   632 => (x"4c",x"a3",x"d0",x"87"),
   633 => (x"bf",x"d2",x"f0",x"c2"),
   634 => (x"6c",x"b9",x"ff",x"49"),
   635 => (x"d4",x"7e",x"99",x"4a"),
   636 => (x"cd",x"06",x"a9",x"66"),
   637 => (x"7c",x"7b",x"c0",x"87"),
   638 => (x"c4",x"4a",x"a3",x"cc"),
   639 => (x"79",x"6a",x"49",x"a3"),
   640 => (x"49",x"72",x"87",x"ca"),
   641 => (x"d4",x"99",x"c0",x"f8"),
   642 => (x"8d",x"71",x"4d",x"66"),
   643 => (x"29",x"c9",x"49",x"75"),
   644 => (x"49",x"73",x"1e",x"71"),
   645 => (x"c2",x"87",x"fa",x"fa"),
   646 => (x"73",x"1e",x"ce",x"e8"),
   647 => (x"87",x"cb",x"fc",x"49"),
   648 => (x"66",x"d4",x"86",x"c8"),
   649 => (x"d6",x"f5",x"26",x"7c"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"c2",x"87",x"e4",x"c0"),
   653 => (x"73",x"5b",x"fb",x"f4"),
   654 => (x"c2",x"8a",x"c2",x"4a"),
   655 => (x"49",x"bf",x"ce",x"f0"),
   656 => (x"e7",x"f4",x"c2",x"92"),
   657 => (x"80",x"72",x"48",x"bf"),
   658 => (x"58",x"ff",x"f4",x"c2"),
   659 => (x"30",x"c4",x"48",x"71"),
   660 => (x"58",x"de",x"f0",x"c2"),
   661 => (x"c2",x"87",x"ed",x"c0"),
   662 => (x"c2",x"48",x"f7",x"f4"),
   663 => (x"78",x"bf",x"eb",x"f4"),
   664 => (x"48",x"fb",x"f4",x"c2"),
   665 => (x"bf",x"ef",x"f4",x"c2"),
   666 => (x"d6",x"f0",x"c2",x"78"),
   667 => (x"87",x"c9",x"02",x"bf"),
   668 => (x"bf",x"ce",x"f0",x"c2"),
   669 => (x"c7",x"31",x"c4",x"49"),
   670 => (x"f3",x"f4",x"c2",x"87"),
   671 => (x"31",x"c4",x"49",x"bf"),
   672 => (x"59",x"de",x"f0",x"c2"),
   673 => (x"0e",x"87",x"fc",x"f3"),
   674 => (x"0e",x"5c",x"5b",x"5e"),
   675 => (x"4b",x"c0",x"4a",x"71"),
   676 => (x"c0",x"02",x"9a",x"72"),
   677 => (x"a2",x"da",x"87",x"e0"),
   678 => (x"4b",x"69",x"9f",x"49"),
   679 => (x"bf",x"d6",x"f0",x"c2"),
   680 => (x"d4",x"87",x"cf",x"02"),
   681 => (x"69",x"9f",x"49",x"a2"),
   682 => (x"ff",x"c0",x"4c",x"49"),
   683 => (x"34",x"d0",x"9c",x"ff"),
   684 => (x"4c",x"c0",x"87",x"c2"),
   685 => (x"49",x"73",x"b3",x"74"),
   686 => (x"f3",x"87",x"ee",x"fd"),
   687 => (x"5e",x"0e",x"87",x"c3"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"4a",x"71",x"86",x"f4"),
   690 => (x"9a",x"72",x"7e",x"c0"),
   691 => (x"c2",x"87",x"d8",x"02"),
   692 => (x"c0",x"48",x"ca",x"e8"),
   693 => (x"c2",x"e8",x"c2",x"78"),
   694 => (x"fb",x"f4",x"c2",x"48"),
   695 => (x"e8",x"c2",x"78",x"bf"),
   696 => (x"f4",x"c2",x"48",x"c6"),
   697 => (x"c2",x"78",x"bf",x"f7"),
   698 => (x"c0",x"48",x"eb",x"f0"),
   699 => (x"da",x"f0",x"c2",x"50"),
   700 => (x"e8",x"c2",x"49",x"bf"),
   701 => (x"71",x"4a",x"bf",x"ca"),
   702 => (x"c9",x"c4",x"03",x"aa"),
   703 => (x"cf",x"49",x"72",x"87"),
   704 => (x"e9",x"c0",x"05",x"99"),
   705 => (x"d5",x"f2",x"c0",x"87"),
   706 => (x"c2",x"e8",x"c2",x"48"),
   707 => (x"e8",x"c2",x"78",x"bf"),
   708 => (x"e8",x"c2",x"1e",x"ce"),
   709 => (x"c2",x"49",x"bf",x"c2"),
   710 => (x"c1",x"48",x"c2",x"e8"),
   711 => (x"e3",x"71",x"78",x"a1"),
   712 => (x"86",x"c4",x"87",x"ed"),
   713 => (x"48",x"d1",x"f2",x"c0"),
   714 => (x"78",x"ce",x"e8",x"c2"),
   715 => (x"f2",x"c0",x"87",x"cc"),
   716 => (x"c0",x"48",x"bf",x"d1"),
   717 => (x"f2",x"c0",x"80",x"e0"),
   718 => (x"e8",x"c2",x"58",x"d5"),
   719 => (x"c1",x"48",x"bf",x"ca"),
   720 => (x"ce",x"e8",x"c2",x"80"),
   721 => (x"0c",x"91",x"27",x"58"),
   722 => (x"97",x"bf",x"00",x"00"),
   723 => (x"02",x"9d",x"4d",x"bf"),
   724 => (x"c3",x"87",x"e3",x"c2"),
   725 => (x"c2",x"02",x"ad",x"e5"),
   726 => (x"f2",x"c0",x"87",x"dc"),
   727 => (x"cb",x"4b",x"bf",x"d1"),
   728 => (x"4c",x"11",x"49",x"a3"),
   729 => (x"c1",x"05",x"ac",x"cf"),
   730 => (x"49",x"75",x"87",x"d2"),
   731 => (x"89",x"c1",x"99",x"df"),
   732 => (x"f0",x"c2",x"91",x"cd"),
   733 => (x"a3",x"c1",x"81",x"de"),
   734 => (x"c3",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"c5"),
   737 => (x"4a",x"a3",x"c7",x"51"),
   738 => (x"a3",x"c9",x"51",x"12"),
   739 => (x"ce",x"51",x"12",x"4a"),
   740 => (x"51",x"12",x"4a",x"a3"),
   741 => (x"12",x"4a",x"a3",x"d0"),
   742 => (x"4a",x"a3",x"d2",x"51"),
   743 => (x"a3",x"d4",x"51",x"12"),
   744 => (x"d6",x"51",x"12",x"4a"),
   745 => (x"51",x"12",x"4a",x"a3"),
   746 => (x"12",x"4a",x"a3",x"d8"),
   747 => (x"4a",x"a3",x"dc",x"51"),
   748 => (x"a3",x"de",x"51",x"12"),
   749 => (x"c1",x"51",x"12",x"4a"),
   750 => (x"87",x"fa",x"c0",x"7e"),
   751 => (x"99",x"c8",x"49",x"74"),
   752 => (x"87",x"eb",x"c0",x"05"),
   753 => (x"99",x"d0",x"49",x"74"),
   754 => (x"dc",x"87",x"d1",x"05"),
   755 => (x"cb",x"c0",x"02",x"66"),
   756 => (x"dc",x"49",x"73",x"87"),
   757 => (x"98",x"70",x"0f",x"66"),
   758 => (x"87",x"d3",x"c0",x"02"),
   759 => (x"c6",x"c0",x"05",x"6e"),
   760 => (x"de",x"f0",x"c2",x"87"),
   761 => (x"c0",x"50",x"c0",x"48"),
   762 => (x"48",x"bf",x"d1",x"f2"),
   763 => (x"c2",x"87",x"dd",x"c2"),
   764 => (x"c0",x"48",x"eb",x"f0"),
   765 => (x"f0",x"c2",x"7e",x"50"),
   766 => (x"c2",x"49",x"bf",x"da"),
   767 => (x"4a",x"bf",x"ca",x"e8"),
   768 => (x"fb",x"04",x"aa",x"71"),
   769 => (x"f4",x"c2",x"87",x"f7"),
   770 => (x"c0",x"05",x"bf",x"fb"),
   771 => (x"f0",x"c2",x"87",x"c8"),
   772 => (x"c1",x"02",x"bf",x"d6"),
   773 => (x"e8",x"c2",x"87",x"f4"),
   774 => (x"ed",x"49",x"bf",x"c6"),
   775 => (x"e8",x"c2",x"87",x"e9"),
   776 => (x"a6",x"c4",x"58",x"ca"),
   777 => (x"c6",x"e8",x"c2",x"48"),
   778 => (x"f0",x"c2",x"78",x"bf"),
   779 => (x"c0",x"02",x"bf",x"d6"),
   780 => (x"66",x"c4",x"87",x"d8"),
   781 => (x"ff",x"ff",x"cf",x"49"),
   782 => (x"a9",x"99",x"f8",x"ff"),
   783 => (x"87",x"c5",x"c0",x"02"),
   784 => (x"e1",x"c0",x"4c",x"c0"),
   785 => (x"c0",x"4c",x"c1",x"87"),
   786 => (x"66",x"c4",x"87",x"dc"),
   787 => (x"f8",x"ff",x"cf",x"49"),
   788 => (x"c0",x"02",x"a9",x"99"),
   789 => (x"a6",x"c8",x"87",x"c8"),
   790 => (x"c0",x"78",x"c0",x"48"),
   791 => (x"a6",x"c8",x"87",x"c5"),
   792 => (x"c8",x"78",x"c1",x"48"),
   793 => (x"9c",x"74",x"4c",x"66"),
   794 => (x"87",x"de",x"c0",x"05"),
   795 => (x"c2",x"49",x"66",x"c4"),
   796 => (x"ce",x"f0",x"c2",x"89"),
   797 => (x"f4",x"c2",x"91",x"bf"),
   798 => (x"71",x"48",x"bf",x"e7"),
   799 => (x"c6",x"e8",x"c2",x"80"),
   800 => (x"ca",x"e8",x"c2",x"58"),
   801 => (x"f9",x"78",x"c0",x"48"),
   802 => (x"48",x"c0",x"87",x"e3"),
   803 => (x"ee",x"eb",x"8e",x"f4"),
   804 => (x"00",x"00",x"00",x"87"),
   805 => (x"ff",x"ff",x"ff",x"00"),
   806 => (x"00",x"0c",x"a1",x"ff"),
   807 => (x"00",x"0c",x"aa",x"00"),
   808 => (x"54",x"41",x"46",x"00"),
   809 => (x"20",x"20",x"32",x"33"),
   810 => (x"41",x"46",x"00",x"20"),
   811 => (x"20",x"36",x"31",x"54"),
   812 => (x"1e",x"00",x"20",x"20"),
   813 => (x"c3",x"48",x"d4",x"ff"),
   814 => (x"48",x"68",x"78",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"ff",x"c3",x"48",x"d4"),
   817 => (x"48",x"d0",x"ff",x"78"),
   818 => (x"ff",x"78",x"e1",x"c0"),
   819 => (x"78",x"d4",x"48",x"d4"),
   820 => (x"48",x"ff",x"f4",x"c2"),
   821 => (x"50",x"bf",x"d4",x"ff"),
   822 => (x"ff",x"1e",x"4f",x"26"),
   823 => (x"e0",x"c0",x"48",x"d0"),
   824 => (x"1e",x"4f",x"26",x"78"),
   825 => (x"70",x"87",x"cc",x"ff"),
   826 => (x"c6",x"02",x"99",x"49"),
   827 => (x"a9",x"fb",x"c0",x"87"),
   828 => (x"71",x"87",x"f1",x"05"),
   829 => (x"0e",x"4f",x"26",x"48"),
   830 => (x"0e",x"5c",x"5b",x"5e"),
   831 => (x"4c",x"c0",x"4b",x"71"),
   832 => (x"70",x"87",x"f0",x"fe"),
   833 => (x"c0",x"02",x"99",x"49"),
   834 => (x"ec",x"c0",x"87",x"f9"),
   835 => (x"f2",x"c0",x"02",x"a9"),
   836 => (x"a9",x"fb",x"c0",x"87"),
   837 => (x"87",x"eb",x"c0",x"02"),
   838 => (x"ac",x"b7",x"66",x"cc"),
   839 => (x"d0",x"87",x"c7",x"03"),
   840 => (x"87",x"c2",x"02",x"66"),
   841 => (x"99",x"71",x"53",x"71"),
   842 => (x"c1",x"87",x"c2",x"02"),
   843 => (x"87",x"c3",x"fe",x"84"),
   844 => (x"02",x"99",x"49",x"70"),
   845 => (x"ec",x"c0",x"87",x"cd"),
   846 => (x"87",x"c7",x"02",x"a9"),
   847 => (x"05",x"a9",x"fb",x"c0"),
   848 => (x"d0",x"87",x"d5",x"ff"),
   849 => (x"87",x"c3",x"02",x"66"),
   850 => (x"c0",x"7b",x"97",x"c0"),
   851 => (x"c4",x"05",x"a9",x"ec"),
   852 => (x"c5",x"4a",x"74",x"87"),
   853 => (x"c0",x"4a",x"74",x"87"),
   854 => (x"48",x"72",x"8a",x"0a"),
   855 => (x"4d",x"26",x"87",x"c2"),
   856 => (x"4b",x"26",x"4c",x"26"),
   857 => (x"fd",x"1e",x"4f",x"26"),
   858 => (x"49",x"70",x"87",x"c9"),
   859 => (x"aa",x"f0",x"c0",x"4a"),
   860 => (x"c0",x"87",x"c9",x"04"),
   861 => (x"c3",x"01",x"aa",x"f9"),
   862 => (x"8a",x"f0",x"c0",x"87"),
   863 => (x"04",x"aa",x"c1",x"c1"),
   864 => (x"da",x"c1",x"87",x"c9"),
   865 => (x"87",x"c3",x"01",x"aa"),
   866 => (x"72",x"8a",x"f7",x"c0"),
   867 => (x"0e",x"4f",x"26",x"48"),
   868 => (x"5d",x"5c",x"5b",x"5e"),
   869 => (x"71",x"86",x"f8",x"0e"),
   870 => (x"c0",x"4d",x"c0",x"4b"),
   871 => (x"bf",x"97",x"e8",x"f9"),
   872 => (x"05",x"a9",x"df",x"49"),
   873 => (x"c8",x"87",x"ee",x"c0"),
   874 => (x"69",x"97",x"49",x"a3"),
   875 => (x"a9",x"c3",x"c1",x"49"),
   876 => (x"c9",x"87",x"dd",x"05"),
   877 => (x"69",x"97",x"49",x"a3"),
   878 => (x"a9",x"c6",x"c1",x"49"),
   879 => (x"ca",x"87",x"d1",x"05"),
   880 => (x"69",x"97",x"49",x"a3"),
   881 => (x"a9",x"c7",x"c1",x"49"),
   882 => (x"c1",x"87",x"c5",x"05"),
   883 => (x"87",x"d3",x"c2",x"48"),
   884 => (x"ce",x"c2",x"48",x"c0"),
   885 => (x"87",x"e6",x"fb",x"87"),
   886 => (x"f9",x"c0",x"4c",x"c0"),
   887 => (x"49",x"bf",x"97",x"e8"),
   888 => (x"cf",x"04",x"a9",x"c0"),
   889 => (x"87",x"fb",x"fb",x"87"),
   890 => (x"f9",x"c0",x"84",x"c1"),
   891 => (x"49",x"bf",x"97",x"e8"),
   892 => (x"87",x"f1",x"06",x"ac"),
   893 => (x"97",x"e8",x"f9",x"c0"),
   894 => (x"87",x"cf",x"02",x"bf"),
   895 => (x"70",x"87",x"f4",x"fa"),
   896 => (x"c6",x"02",x"99",x"49"),
   897 => (x"a9",x"ec",x"c0",x"87"),
   898 => (x"c0",x"87",x"f1",x"05"),
   899 => (x"87",x"e3",x"fa",x"4c"),
   900 => (x"de",x"fa",x"7e",x"70"),
   901 => (x"58",x"a6",x"c8",x"87"),
   902 => (x"70",x"87",x"d8",x"fa"),
   903 => (x"c8",x"84",x"c1",x"4a"),
   904 => (x"69",x"97",x"49",x"a3"),
   905 => (x"05",x"a9",x"6e",x"49"),
   906 => (x"a3",x"c9",x"87",x"da"),
   907 => (x"49",x"69",x"97",x"49"),
   908 => (x"05",x"a9",x"66",x"c4"),
   909 => (x"a3",x"ca",x"87",x"ce"),
   910 => (x"49",x"69",x"97",x"49"),
   911 => (x"87",x"c4",x"05",x"aa"),
   912 => (x"87",x"d4",x"4d",x"c1"),
   913 => (x"ec",x"c0",x"48",x"6e"),
   914 => (x"87",x"c8",x"02",x"a8"),
   915 => (x"fb",x"c0",x"48",x"6e"),
   916 => (x"87",x"c4",x"05",x"a8"),
   917 => (x"4d",x"c1",x"4c",x"c0"),
   918 => (x"fe",x"02",x"9d",x"75"),
   919 => (x"f9",x"f9",x"87",x"ef"),
   920 => (x"f8",x"48",x"74",x"87"),
   921 => (x"87",x"f6",x"fb",x"8e"),
   922 => (x"5b",x"5e",x"0e",x"00"),
   923 => (x"f8",x"0e",x"5d",x"5c"),
   924 => (x"ff",x"7e",x"71",x"86"),
   925 => (x"1e",x"6e",x"4b",x"d4"),
   926 => (x"49",x"c4",x"f5",x"c2"),
   927 => (x"c4",x"87",x"fa",x"e5"),
   928 => (x"02",x"98",x"70",x"86"),
   929 => (x"c1",x"87",x"ea",x"c4"),
   930 => (x"4d",x"bf",x"ce",x"e7"),
   931 => (x"fe",x"fb",x"49",x"6e"),
   932 => (x"58",x"a6",x"c8",x"87"),
   933 => (x"c5",x"05",x"98",x"70"),
   934 => (x"48",x"a6",x"c4",x"87"),
   935 => (x"d0",x"ff",x"78",x"c1"),
   936 => (x"c1",x"78",x"c5",x"48"),
   937 => (x"66",x"c4",x"7b",x"d5"),
   938 => (x"c6",x"89",x"c1",x"49"),
   939 => (x"cc",x"e7",x"c1",x"31"),
   940 => (x"48",x"4a",x"bf",x"97"),
   941 => (x"7b",x"70",x"b0",x"71"),
   942 => (x"c4",x"48",x"d0",x"ff"),
   943 => (x"ff",x"f4",x"c2",x"78"),
   944 => (x"d0",x"49",x"bf",x"97"),
   945 => (x"87",x"d7",x"02",x"99"),
   946 => (x"d6",x"c1",x"78",x"c5"),
   947 => (x"c3",x"4a",x"c0",x"7b"),
   948 => (x"82",x"c1",x"7b",x"ff"),
   949 => (x"04",x"aa",x"e0",x"c0"),
   950 => (x"d0",x"ff",x"87",x"f5"),
   951 => (x"c3",x"78",x"c4",x"48"),
   952 => (x"d0",x"ff",x"7b",x"ff"),
   953 => (x"c1",x"78",x"c5",x"48"),
   954 => (x"7b",x"c1",x"7b",x"d3"),
   955 => (x"b7",x"c0",x"78",x"c4"),
   956 => (x"eb",x"c2",x"06",x"ad"),
   957 => (x"cc",x"f5",x"c2",x"87"),
   958 => (x"9c",x"8d",x"4c",x"bf"),
   959 => (x"87",x"c2",x"c2",x"02"),
   960 => (x"7e",x"ce",x"e8",x"c2"),
   961 => (x"c8",x"48",x"a6",x"c4"),
   962 => (x"c0",x"8c",x"78",x"c0"),
   963 => (x"c6",x"03",x"ac",x"b7"),
   964 => (x"a4",x"c0",x"c8",x"87"),
   965 => (x"c2",x"4c",x"c0",x"78"),
   966 => (x"bf",x"97",x"ff",x"f4"),
   967 => (x"02",x"99",x"d0",x"49"),
   968 => (x"1e",x"c0",x"87",x"d0"),
   969 => (x"49",x"c4",x"f5",x"c2"),
   970 => (x"c4",x"87",x"c0",x"e8"),
   971 => (x"c0",x"4a",x"70",x"86"),
   972 => (x"e8",x"c2",x"87",x"f5"),
   973 => (x"f5",x"c2",x"1e",x"ce"),
   974 => (x"ee",x"e7",x"49",x"c4"),
   975 => (x"70",x"86",x"c4",x"87"),
   976 => (x"48",x"d0",x"ff",x"4a"),
   977 => (x"c1",x"78",x"c5",x"c8"),
   978 => (x"97",x"6e",x"7b",x"d4"),
   979 => (x"48",x"6e",x"7b",x"bf"),
   980 => (x"7e",x"70",x"80",x"c1"),
   981 => (x"c1",x"48",x"66",x"c4"),
   982 => (x"58",x"a6",x"c8",x"88"),
   983 => (x"ff",x"05",x"98",x"70"),
   984 => (x"d0",x"ff",x"87",x"e8"),
   985 => (x"72",x"78",x"c4",x"48"),
   986 => (x"87",x"c5",x"05",x"9a"),
   987 => (x"c2",x"c1",x"48",x"c0"),
   988 => (x"c2",x"1e",x"c1",x"87"),
   989 => (x"e5",x"49",x"c4",x"f5"),
   990 => (x"86",x"c4",x"87",x"d7"),
   991 => (x"fd",x"05",x"9c",x"74"),
   992 => (x"b7",x"c0",x"87",x"fe"),
   993 => (x"87",x"d1",x"06",x"ad"),
   994 => (x"48",x"c4",x"f5",x"c2"),
   995 => (x"80",x"d0",x"78",x"c0"),
   996 => (x"80",x"f4",x"78",x"c0"),
   997 => (x"bf",x"d0",x"f5",x"c2"),
   998 => (x"ad",x"b7",x"c0",x"78"),
   999 => (x"87",x"d5",x"fd",x"01"),
  1000 => (x"c5",x"48",x"d0",x"ff"),
  1001 => (x"7b",x"d3",x"c1",x"78"),
  1002 => (x"78",x"c4",x"7b",x"c0"),
  1003 => (x"c2",x"c0",x"48",x"c1"),
  1004 => (x"f8",x"48",x"c0",x"87"),
  1005 => (x"26",x"4d",x"26",x"8e"),
  1006 => (x"26",x"4b",x"26",x"4c"),
  1007 => (x"5b",x"5e",x"0e",x"4f"),
  1008 => (x"1e",x"0e",x"5d",x"5c"),
  1009 => (x"4c",x"c0",x"4b",x"71"),
  1010 => (x"c0",x"04",x"ab",x"4d"),
  1011 => (x"f6",x"c0",x"87",x"e8"),
  1012 => (x"9d",x"75",x"1e",x"cf"),
  1013 => (x"c0",x"87",x"c4",x"02"),
  1014 => (x"c1",x"87",x"c2",x"4a"),
  1015 => (x"eb",x"49",x"72",x"4a"),
  1016 => (x"86",x"c4",x"87",x"dc"),
  1017 => (x"84",x"c1",x"7e",x"70"),
  1018 => (x"87",x"c2",x"05",x"6e"),
  1019 => (x"85",x"c1",x"4c",x"73"),
  1020 => (x"ff",x"06",x"ac",x"73"),
  1021 => (x"48",x"6e",x"87",x"d8"),
  1022 => (x"87",x"f9",x"fe",x"26"),
  1023 => (x"5c",x"5b",x"5e",x"0e"),
  1024 => (x"cc",x"4b",x"71",x"0e"),
  1025 => (x"e8",x"c0",x"02",x"66"),
  1026 => (x"f0",x"c0",x"4c",x"87"),
  1027 => (x"e8",x"c0",x"02",x"8c"),
  1028 => (x"c1",x"4a",x"74",x"87"),
  1029 => (x"e0",x"c0",x"02",x"8a"),
  1030 => (x"dc",x"02",x"8a",x"87"),
  1031 => (x"d8",x"02",x"8a",x"87"),
  1032 => (x"8a",x"e0",x"c0",x"87"),
  1033 => (x"87",x"e5",x"c0",x"02"),
  1034 => (x"c0",x"02",x"8a",x"c1"),
  1035 => (x"ea",x"c0",x"87",x"e7"),
  1036 => (x"f8",x"49",x"73",x"87"),
  1037 => (x"e2",x"c0",x"87",x"f3"),
  1038 => (x"c0",x"1e",x"74",x"87"),
  1039 => (x"ce",x"de",x"c1",x"49"),
  1040 => (x"73",x"1e",x"74",x"87"),
  1041 => (x"c6",x"de",x"c1",x"49"),
  1042 => (x"ce",x"86",x"c8",x"87"),
  1043 => (x"c1",x"49",x"73",x"87"),
  1044 => (x"c6",x"87",x"eb",x"e0"),
  1045 => (x"c1",x"49",x"73",x"87"),
  1046 => (x"fd",x"87",x"dd",x"e1"),
  1047 => (x"5e",x"0e",x"87",x"d9"),
  1048 => (x"0e",x"5d",x"5c",x"5b"),
  1049 => (x"49",x"4c",x"71",x"1e"),
  1050 => (x"f5",x"c2",x"91",x"de"),
  1051 => (x"85",x"71",x"4d",x"ec"),
  1052 => (x"c1",x"02",x"6d",x"97"),
  1053 => (x"f5",x"c2",x"87",x"dd"),
  1054 => (x"74",x"49",x"bf",x"d8"),
  1055 => (x"fc",x"fc",x"71",x"81"),
  1056 => (x"48",x"7e",x"70",x"87"),
  1057 => (x"f2",x"c0",x"02",x"98"),
  1058 => (x"e0",x"f5",x"c2",x"87"),
  1059 => (x"cb",x"4a",x"70",x"4b"),
  1060 => (x"d2",x"c0",x"ff",x"49"),
  1061 => (x"cb",x"4b",x"74",x"87"),
  1062 => (x"c3",x"e8",x"c1",x"93"),
  1063 => (x"c1",x"83",x"c4",x"83"),
  1064 => (x"74",x"7b",x"d7",x"c3"),
  1065 => (x"fe",x"c2",x"c1",x"49"),
  1066 => (x"c1",x"7b",x"75",x"87"),
  1067 => (x"bf",x"97",x"cd",x"e7"),
  1068 => (x"f5",x"c2",x"1e",x"49"),
  1069 => (x"c3",x"fd",x"49",x"e0"),
  1070 => (x"74",x"86",x"c4",x"87"),
  1071 => (x"e6",x"c2",x"c1",x"49"),
  1072 => (x"c1",x"49",x"c0",x"87"),
  1073 => (x"c2",x"87",x"c5",x"c4"),
  1074 => (x"c0",x"48",x"c0",x"f5"),
  1075 => (x"c0",x"49",x"c1",x"78"),
  1076 => (x"26",x"87",x"e5",x"e0"),
  1077 => (x"4c",x"87",x"de",x"fb"),
  1078 => (x"69",x"64",x"61",x"6f"),
  1079 => (x"2e",x"2e",x"67",x"6e"),
  1080 => (x"73",x"1e",x"00",x"2e"),
  1081 => (x"49",x"4a",x"71",x"1e"),
  1082 => (x"bf",x"d8",x"f5",x"c2"),
  1083 => (x"cc",x"fb",x"71",x"81"),
  1084 => (x"9b",x"4b",x"70",x"87"),
  1085 => (x"49",x"87",x"c4",x"02"),
  1086 => (x"c2",x"87",x"cc",x"e6"),
  1087 => (x"c0",x"48",x"d8",x"f5"),
  1088 => (x"df",x"49",x"c1",x"78"),
  1089 => (x"f0",x"fa",x"87",x"f2"),
  1090 => (x"49",x"c0",x"1e",x"87"),
  1091 => (x"87",x"fc",x"c2",x"c1"),
  1092 => (x"71",x"1e",x"4f",x"26"),
  1093 => (x"91",x"cb",x"49",x"4a"),
  1094 => (x"81",x"c3",x"e8",x"c1"),
  1095 => (x"48",x"11",x"81",x"c8"),
  1096 => (x"58",x"c4",x"f5",x"c2"),
  1097 => (x"48",x"d8",x"f5",x"c2"),
  1098 => (x"49",x"c1",x"78",x"c0"),
  1099 => (x"26",x"87",x"c9",x"df"),
  1100 => (x"99",x"71",x"1e",x"4f"),
  1101 => (x"c1",x"87",x"d2",x"02"),
  1102 => (x"c0",x"48",x"d8",x"e9"),
  1103 => (x"c1",x"80",x"f7",x"50"),
  1104 => (x"c1",x"40",x"d2",x"c4"),
  1105 => (x"ce",x"78",x"f1",x"e7"),
  1106 => (x"d4",x"e9",x"c1",x"87"),
  1107 => (x"d2",x"e7",x"c1",x"48"),
  1108 => (x"c1",x"80",x"fc",x"78"),
  1109 => (x"26",x"78",x"c9",x"c4"),
  1110 => (x"5b",x"5e",x"0e",x"4f"),
  1111 => (x"f4",x"0e",x"5d",x"5c"),
  1112 => (x"ce",x"e8",x"c2",x"86"),
  1113 => (x"c4",x"4c",x"c0",x"4d"),
  1114 => (x"78",x"c0",x"48",x"a6"),
  1115 => (x"bf",x"d8",x"f5",x"c2"),
  1116 => (x"06",x"a8",x"c0",x"48"),
  1117 => (x"c2",x"87",x"c0",x"c1"),
  1118 => (x"98",x"48",x"ce",x"e8"),
  1119 => (x"87",x"f7",x"c0",x"02"),
  1120 => (x"1e",x"cf",x"f6",x"c0"),
  1121 => (x"c7",x"02",x"66",x"c8"),
  1122 => (x"48",x"a6",x"c4",x"87"),
  1123 => (x"87",x"c5",x"78",x"c0"),
  1124 => (x"c1",x"48",x"a6",x"c4"),
  1125 => (x"49",x"66",x"c4",x"78"),
  1126 => (x"c4",x"87",x"e3",x"e4"),
  1127 => (x"c1",x"4d",x"70",x"86"),
  1128 => (x"48",x"66",x"c4",x"84"),
  1129 => (x"a6",x"c8",x"80",x"c1"),
  1130 => (x"d8",x"f5",x"c2",x"58"),
  1131 => (x"c6",x"03",x"ac",x"bf"),
  1132 => (x"05",x"9d",x"75",x"87"),
  1133 => (x"c0",x"87",x"c9",x"ff"),
  1134 => (x"02",x"9d",x"75",x"4c"),
  1135 => (x"c0",x"87",x"dc",x"c3"),
  1136 => (x"c8",x"1e",x"cf",x"f6"),
  1137 => (x"87",x"c7",x"02",x"66"),
  1138 => (x"c0",x"48",x"a6",x"cc"),
  1139 => (x"cc",x"87",x"c5",x"78"),
  1140 => (x"78",x"c1",x"48",x"a6"),
  1141 => (x"e3",x"49",x"66",x"cc"),
  1142 => (x"86",x"c4",x"87",x"e4"),
  1143 => (x"98",x"48",x"7e",x"70"),
  1144 => (x"87",x"e4",x"c2",x"02"),
  1145 => (x"97",x"81",x"cb",x"49"),
  1146 => (x"99",x"d0",x"49",x"69"),
  1147 => (x"87",x"d4",x"c1",x"02"),
  1148 => (x"91",x"cb",x"49",x"74"),
  1149 => (x"81",x"c3",x"e8",x"c1"),
  1150 => (x"79",x"e2",x"c3",x"c1"),
  1151 => (x"ff",x"c3",x"81",x"c8"),
  1152 => (x"de",x"49",x"74",x"51"),
  1153 => (x"ec",x"f5",x"c2",x"91"),
  1154 => (x"c2",x"85",x"71",x"4d"),
  1155 => (x"c1",x"7d",x"97",x"c1"),
  1156 => (x"e0",x"c0",x"49",x"a5"),
  1157 => (x"de",x"f0",x"c2",x"51"),
  1158 => (x"d2",x"02",x"bf",x"97"),
  1159 => (x"c2",x"84",x"c1",x"87"),
  1160 => (x"f0",x"c2",x"4b",x"a5"),
  1161 => (x"49",x"db",x"4a",x"de"),
  1162 => (x"87",x"fb",x"f9",x"fe"),
  1163 => (x"cd",x"87",x"d9",x"c1"),
  1164 => (x"51",x"c0",x"49",x"a5"),
  1165 => (x"a5",x"c2",x"84",x"c1"),
  1166 => (x"cb",x"4a",x"6e",x"4b"),
  1167 => (x"e6",x"f9",x"fe",x"49"),
  1168 => (x"87",x"c4",x"c1",x"87"),
  1169 => (x"91",x"cb",x"49",x"74"),
  1170 => (x"81",x"c3",x"e8",x"c1"),
  1171 => (x"79",x"de",x"c1",x"c1"),
  1172 => (x"97",x"de",x"f0",x"c2"),
  1173 => (x"87",x"d8",x"02",x"bf"),
  1174 => (x"91",x"de",x"49",x"74"),
  1175 => (x"f5",x"c2",x"84",x"c1"),
  1176 => (x"83",x"71",x"4b",x"ec"),
  1177 => (x"4a",x"de",x"f0",x"c2"),
  1178 => (x"f8",x"fe",x"49",x"dd"),
  1179 => (x"87",x"d8",x"87",x"f9"),
  1180 => (x"93",x"de",x"4b",x"74"),
  1181 => (x"83",x"ec",x"f5",x"c2"),
  1182 => (x"c0",x"49",x"a3",x"cb"),
  1183 => (x"73",x"84",x"c1",x"51"),
  1184 => (x"49",x"cb",x"4a",x"6e"),
  1185 => (x"87",x"df",x"f8",x"fe"),
  1186 => (x"c1",x"48",x"66",x"c4"),
  1187 => (x"58",x"a6",x"c8",x"80"),
  1188 => (x"c0",x"03",x"ac",x"c7"),
  1189 => (x"05",x"6e",x"87",x"c5"),
  1190 => (x"74",x"87",x"e4",x"fc"),
  1191 => (x"f4",x"8e",x"f4",x"48"),
  1192 => (x"73",x"1e",x"87",x"d3"),
  1193 => (x"49",x"4b",x"71",x"1e"),
  1194 => (x"e8",x"c1",x"91",x"cb"),
  1195 => (x"a1",x"c8",x"81",x"c3"),
  1196 => (x"cc",x"e7",x"c1",x"4a"),
  1197 => (x"c9",x"50",x"12",x"48"),
  1198 => (x"f9",x"c0",x"4a",x"a1"),
  1199 => (x"50",x"12",x"48",x"e8"),
  1200 => (x"e7",x"c1",x"81",x"ca"),
  1201 => (x"50",x"11",x"48",x"cd"),
  1202 => (x"97",x"cd",x"e7",x"c1"),
  1203 => (x"c0",x"1e",x"49",x"bf"),
  1204 => (x"87",x"e8",x"f4",x"49"),
  1205 => (x"48",x"c0",x"f5",x"c2"),
  1206 => (x"49",x"c1",x"78",x"de"),
  1207 => (x"26",x"87",x"d9",x"d8"),
  1208 => (x"0e",x"87",x"d6",x"f3"),
  1209 => (x"5d",x"5c",x"5b",x"5e"),
  1210 => (x"71",x"86",x"f4",x"0e"),
  1211 => (x"91",x"cb",x"49",x"4d"),
  1212 => (x"81",x"c3",x"e8",x"c1"),
  1213 => (x"ca",x"4a",x"a1",x"c8"),
  1214 => (x"a6",x"c4",x"7e",x"a1"),
  1215 => (x"c8",x"f9",x"c2",x"48"),
  1216 => (x"97",x"6e",x"78",x"bf"),
  1217 => (x"66",x"c4",x"4b",x"bf"),
  1218 => (x"12",x"2c",x"73",x"4c"),
  1219 => (x"58",x"a6",x"cc",x"48"),
  1220 => (x"84",x"c1",x"9c",x"70"),
  1221 => (x"69",x"97",x"81",x"c9"),
  1222 => (x"04",x"ac",x"b7",x"49"),
  1223 => (x"4c",x"c0",x"87",x"c2"),
  1224 => (x"4a",x"bf",x"97",x"6e"),
  1225 => (x"72",x"49",x"66",x"c8"),
  1226 => (x"c4",x"b9",x"ff",x"31"),
  1227 => (x"48",x"74",x"99",x"66"),
  1228 => (x"4a",x"70",x"30",x"72"),
  1229 => (x"c2",x"b0",x"71",x"48"),
  1230 => (x"c0",x"58",x"cc",x"f9"),
  1231 => (x"c0",x"87",x"e8",x"e6"),
  1232 => (x"87",x"f4",x"d6",x"49"),
  1233 => (x"f8",x"c0",x"49",x"75"),
  1234 => (x"8e",x"f4",x"87",x"dd"),
  1235 => (x"1e",x"87",x"e6",x"f1"),
  1236 => (x"4b",x"71",x"1e",x"73"),
  1237 => (x"87",x"cb",x"fe",x"49"),
  1238 => (x"c6",x"fe",x"49",x"73"),
  1239 => (x"87",x"d9",x"f1",x"87"),
  1240 => (x"71",x"1e",x"73",x"1e"),
  1241 => (x"4a",x"a3",x"c6",x"4b"),
  1242 => (x"87",x"e3",x"c0",x"02"),
  1243 => (x"d6",x"02",x"8a",x"c1"),
  1244 => (x"c1",x"02",x"8a",x"87"),
  1245 => (x"02",x"8a",x"87",x"e8"),
  1246 => (x"8a",x"87",x"ca",x"c1"),
  1247 => (x"87",x"ef",x"c0",x"02"),
  1248 => (x"87",x"d9",x"02",x"8a"),
  1249 => (x"c7",x"87",x"e9",x"c1"),
  1250 => (x"87",x"c6",x"f6",x"49"),
  1251 => (x"c2",x"87",x"ec",x"c1"),
  1252 => (x"df",x"48",x"c0",x"f5"),
  1253 => (x"d5",x"49",x"c1",x"78"),
  1254 => (x"de",x"c1",x"87",x"de"),
  1255 => (x"d8",x"f5",x"c2",x"87"),
  1256 => (x"cb",x"c1",x"02",x"bf"),
  1257 => (x"88",x"c1",x"48",x"87"),
  1258 => (x"58",x"dc",x"f5",x"c2"),
  1259 => (x"c2",x"87",x"c1",x"c1"),
  1260 => (x"02",x"bf",x"dc",x"f5"),
  1261 => (x"c2",x"87",x"f9",x"c0"),
  1262 => (x"48",x"bf",x"d8",x"f5"),
  1263 => (x"f5",x"c2",x"80",x"c1"),
  1264 => (x"eb",x"c0",x"58",x"dc"),
  1265 => (x"d8",x"f5",x"c2",x"87"),
  1266 => (x"89",x"c6",x"49",x"bf"),
  1267 => (x"59",x"dc",x"f5",x"c2"),
  1268 => (x"03",x"a9",x"b7",x"c0"),
  1269 => (x"f5",x"c2",x"87",x"da"),
  1270 => (x"78",x"c0",x"48",x"d8"),
  1271 => (x"f5",x"c2",x"87",x"d2"),
  1272 => (x"cb",x"02",x"bf",x"dc"),
  1273 => (x"d8",x"f5",x"c2",x"87"),
  1274 => (x"80",x"c6",x"48",x"bf"),
  1275 => (x"58",x"dc",x"f5",x"c2"),
  1276 => (x"c3",x"d4",x"49",x"c0"),
  1277 => (x"c0",x"49",x"73",x"87"),
  1278 => (x"ee",x"87",x"ec",x"f5"),
  1279 => (x"5e",x"0e",x"87",x"fb"),
  1280 => (x"0e",x"5d",x"5c",x"5b"),
  1281 => (x"dc",x"86",x"d4",x"ff"),
  1282 => (x"a6",x"c8",x"59",x"a6"),
  1283 => (x"c4",x"78",x"c0",x"48"),
  1284 => (x"66",x"c0",x"c1",x"80"),
  1285 => (x"c1",x"80",x"c4",x"78"),
  1286 => (x"c1",x"80",x"c4",x"78"),
  1287 => (x"dc",x"f5",x"c2",x"78"),
  1288 => (x"c2",x"78",x"c1",x"48"),
  1289 => (x"7e",x"bf",x"c0",x"f5"),
  1290 => (x"a8",x"de",x"48",x"6e"),
  1291 => (x"f4",x"87",x"c9",x"05"),
  1292 => (x"a6",x"cc",x"87",x"e7"),
  1293 => (x"87",x"df",x"d1",x"58"),
  1294 => (x"a8",x"df",x"48",x"6e"),
  1295 => (x"87",x"ea",x"c1",x"05"),
  1296 => (x"49",x"66",x"fc",x"c0"),
  1297 => (x"7e",x"69",x"81",x"c4"),
  1298 => (x"48",x"cc",x"e3",x"c1"),
  1299 => (x"a1",x"d0",x"49",x"6e"),
  1300 => (x"71",x"41",x"20",x"4a"),
  1301 => (x"87",x"f9",x"05",x"aa"),
  1302 => (x"48",x"66",x"fc",x"c0"),
  1303 => (x"78",x"e2",x"ca",x"c1"),
  1304 => (x"49",x"66",x"fc",x"c0"),
  1305 => (x"51",x"df",x"81",x"c9"),
  1306 => (x"49",x"66",x"fc",x"c0"),
  1307 => (x"d3",x"c1",x"81",x"ca"),
  1308 => (x"66",x"fc",x"c0",x"51"),
  1309 => (x"c4",x"81",x"cb",x"49"),
  1310 => (x"a6",x"c4",x"4a",x"a1"),
  1311 => (x"71",x"78",x"6a",x"48"),
  1312 => (x"dc",x"e3",x"c1",x"1e"),
  1313 => (x"49",x"66",x"c8",x"48"),
  1314 => (x"20",x"4a",x"a1",x"d0"),
  1315 => (x"05",x"aa",x"71",x"41"),
  1316 => (x"49",x"26",x"87",x"f9"),
  1317 => (x"79",x"e2",x"ca",x"c1"),
  1318 => (x"df",x"4a",x"a1",x"c9"),
  1319 => (x"c1",x"81",x"ca",x"52"),
  1320 => (x"a6",x"c8",x"51",x"d4"),
  1321 => (x"cf",x"78",x"c2",x"48"),
  1322 => (x"d1",x"e0",x"87",x"ed"),
  1323 => (x"87",x"f3",x"e0",x"87"),
  1324 => (x"70",x"87",x"c0",x"e0"),
  1325 => (x"ac",x"fb",x"c0",x"4c"),
  1326 => (x"87",x"fd",x"c1",x"02"),
  1327 => (x"c1",x"05",x"66",x"d8"),
  1328 => (x"fc",x"c0",x"87",x"ee"),
  1329 => (x"82",x"c4",x"4a",x"66"),
  1330 => (x"1e",x"72",x"7e",x"6a"),
  1331 => (x"48",x"ec",x"e3",x"c1"),
  1332 => (x"c8",x"49",x"66",x"c4"),
  1333 => (x"41",x"20",x"4a",x"a1"),
  1334 => (x"f9",x"05",x"aa",x"71"),
  1335 => (x"26",x"51",x"10",x"87"),
  1336 => (x"66",x"fc",x"c0",x"4a"),
  1337 => (x"e2",x"ca",x"c1",x"48"),
  1338 => (x"c7",x"49",x"6a",x"78"),
  1339 => (x"c0",x"51",x"74",x"81"),
  1340 => (x"c8",x"49",x"66",x"fc"),
  1341 => (x"c0",x"51",x"c1",x"81"),
  1342 => (x"c9",x"49",x"66",x"fc"),
  1343 => (x"c0",x"51",x"c0",x"81"),
  1344 => (x"ca",x"49",x"66",x"fc"),
  1345 => (x"c1",x"51",x"c0",x"81"),
  1346 => (x"6a",x"1e",x"d8",x"1e"),
  1347 => (x"ff",x"81",x"c8",x"49"),
  1348 => (x"c8",x"87",x"e4",x"df"),
  1349 => (x"66",x"c0",x"c1",x"86"),
  1350 => (x"01",x"a8",x"c0",x"48"),
  1351 => (x"a6",x"c8",x"87",x"c7"),
  1352 => (x"cf",x"78",x"c1",x"48"),
  1353 => (x"66",x"c0",x"c1",x"87"),
  1354 => (x"d0",x"88",x"c1",x"48"),
  1355 => (x"87",x"c4",x"58",x"a6"),
  1356 => (x"87",x"ef",x"de",x"ff"),
  1357 => (x"c2",x"48",x"a6",x"d0"),
  1358 => (x"02",x"9c",x"74",x"78"),
  1359 => (x"c8",x"87",x"d4",x"cd"),
  1360 => (x"c4",x"c1",x"48",x"66"),
  1361 => (x"cd",x"03",x"a8",x"66"),
  1362 => (x"a6",x"dc",x"87",x"c9"),
  1363 => (x"e8",x"78",x"c0",x"48"),
  1364 => (x"ff",x"78",x"c0",x"80"),
  1365 => (x"70",x"87",x"dc",x"dd"),
  1366 => (x"ac",x"d0",x"c1",x"4c"),
  1367 => (x"87",x"d9",x"c2",x"05"),
  1368 => (x"e0",x"7e",x"66",x"c4"),
  1369 => (x"a6",x"c8",x"87",x"c0"),
  1370 => (x"c6",x"dd",x"ff",x"58"),
  1371 => (x"c0",x"4c",x"70",x"87"),
  1372 => (x"c1",x"05",x"ac",x"ec"),
  1373 => (x"66",x"c8",x"87",x"ed"),
  1374 => (x"c0",x"91",x"cb",x"49"),
  1375 => (x"c4",x"81",x"66",x"fc"),
  1376 => (x"4d",x"6a",x"4a",x"a1"),
  1377 => (x"c4",x"4a",x"a1",x"c8"),
  1378 => (x"c4",x"c1",x"52",x"66"),
  1379 => (x"dc",x"ff",x"79",x"d2"),
  1380 => (x"4c",x"70",x"87",x"e1"),
  1381 => (x"87",x"d9",x"02",x"9c"),
  1382 => (x"02",x"ac",x"fb",x"c0"),
  1383 => (x"55",x"74",x"87",x"d3"),
  1384 => (x"87",x"cf",x"dc",x"ff"),
  1385 => (x"02",x"9c",x"4c",x"70"),
  1386 => (x"fb",x"c0",x"87",x"c7"),
  1387 => (x"ed",x"ff",x"05",x"ac"),
  1388 => (x"55",x"e0",x"c0",x"87"),
  1389 => (x"c0",x"55",x"c1",x"c2"),
  1390 => (x"66",x"d8",x"7d",x"97"),
  1391 => (x"05",x"a8",x"6e",x"48"),
  1392 => (x"66",x"c8",x"87",x"db"),
  1393 => (x"a8",x"66",x"cc",x"48"),
  1394 => (x"c8",x"87",x"ca",x"04"),
  1395 => (x"80",x"c1",x"48",x"66"),
  1396 => (x"c8",x"58",x"a6",x"cc"),
  1397 => (x"48",x"66",x"cc",x"87"),
  1398 => (x"a6",x"d0",x"88",x"c1"),
  1399 => (x"d2",x"db",x"ff",x"58"),
  1400 => (x"c1",x"4c",x"70",x"87"),
  1401 => (x"c0",x"05",x"ac",x"d0"),
  1402 => (x"66",x"d4",x"87",x"c8"),
  1403 => (x"d8",x"80",x"c1",x"48"),
  1404 => (x"d0",x"c1",x"58",x"a6"),
  1405 => (x"e7",x"fd",x"02",x"ac"),
  1406 => (x"48",x"66",x"c4",x"87"),
  1407 => (x"05",x"a8",x"66",x"d8"),
  1408 => (x"c0",x"87",x"e2",x"c9"),
  1409 => (x"c0",x"48",x"a6",x"e0"),
  1410 => (x"c0",x"48",x"74",x"78"),
  1411 => (x"7e",x"70",x"88",x"fb"),
  1412 => (x"c9",x"02",x"98",x"48"),
  1413 => (x"cb",x"48",x"87",x"e4"),
  1414 => (x"48",x"7e",x"70",x"88"),
  1415 => (x"cf",x"c1",x"02",x"98"),
  1416 => (x"88",x"c9",x"48",x"87"),
  1417 => (x"98",x"48",x"7e",x"70"),
  1418 => (x"87",x"c0",x"c4",x"02"),
  1419 => (x"70",x"88",x"c4",x"48"),
  1420 => (x"02",x"98",x"48",x"7e"),
  1421 => (x"48",x"87",x"ce",x"c0"),
  1422 => (x"7e",x"70",x"88",x"c1"),
  1423 => (x"c3",x"02",x"98",x"48"),
  1424 => (x"d7",x"c8",x"87",x"ea"),
  1425 => (x"48",x"a6",x"dc",x"87"),
  1426 => (x"ff",x"78",x"f0",x"c0"),
  1427 => (x"70",x"87",x"e4",x"d9"),
  1428 => (x"ac",x"ec",x"c0",x"4c"),
  1429 => (x"87",x"c4",x"c0",x"02"),
  1430 => (x"5c",x"a6",x"e0",x"c0"),
  1431 => (x"02",x"ac",x"ec",x"c0"),
  1432 => (x"ff",x"87",x"cd",x"c0"),
  1433 => (x"70",x"87",x"cc",x"d9"),
  1434 => (x"ac",x"ec",x"c0",x"4c"),
  1435 => (x"87",x"f3",x"ff",x"05"),
  1436 => (x"02",x"ac",x"ec",x"c0"),
  1437 => (x"ff",x"87",x"c4",x"c0"),
  1438 => (x"c0",x"87",x"f8",x"d8"),
  1439 => (x"d0",x"1e",x"ca",x"1e"),
  1440 => (x"91",x"cb",x"49",x"66"),
  1441 => (x"48",x"66",x"c4",x"c1"),
  1442 => (x"a6",x"cc",x"80",x"71"),
  1443 => (x"48",x"66",x"c8",x"58"),
  1444 => (x"a6",x"d0",x"80",x"c4"),
  1445 => (x"bf",x"66",x"cc",x"58"),
  1446 => (x"da",x"d9",x"ff",x"49"),
  1447 => (x"de",x"1e",x"c1",x"87"),
  1448 => (x"bf",x"66",x"d4",x"1e"),
  1449 => (x"ce",x"d9",x"ff",x"49"),
  1450 => (x"70",x"86",x"d0",x"87"),
  1451 => (x"08",x"c0",x"48",x"49"),
  1452 => (x"a6",x"e8",x"c0",x"88"),
  1453 => (x"06",x"a8",x"c0",x"58"),
  1454 => (x"c0",x"87",x"ee",x"c0"),
  1455 => (x"dd",x"48",x"66",x"e4"),
  1456 => (x"e4",x"c0",x"03",x"a8"),
  1457 => (x"bf",x"66",x"c4",x"87"),
  1458 => (x"66",x"e4",x"c0",x"49"),
  1459 => (x"51",x"e0",x"c0",x"81"),
  1460 => (x"49",x"66",x"e4",x"c0"),
  1461 => (x"66",x"c4",x"81",x"c1"),
  1462 => (x"c1",x"c2",x"81",x"bf"),
  1463 => (x"66",x"e4",x"c0",x"51"),
  1464 => (x"c4",x"81",x"c2",x"49"),
  1465 => (x"c0",x"81",x"bf",x"66"),
  1466 => (x"c1",x"48",x"6e",x"51"),
  1467 => (x"6e",x"78",x"e2",x"ca"),
  1468 => (x"d0",x"81",x"c8",x"49"),
  1469 => (x"49",x"6e",x"51",x"66"),
  1470 => (x"66",x"d4",x"81",x"c9"),
  1471 => (x"ca",x"49",x"6e",x"51"),
  1472 => (x"51",x"66",x"dc",x"81"),
  1473 => (x"c1",x"48",x"66",x"d0"),
  1474 => (x"58",x"a6",x"d4",x"80"),
  1475 => (x"cc",x"48",x"66",x"c8"),
  1476 => (x"c0",x"04",x"a8",x"66"),
  1477 => (x"66",x"c8",x"87",x"cb"),
  1478 => (x"cc",x"80",x"c1",x"48"),
  1479 => (x"d9",x"c5",x"58",x"a6"),
  1480 => (x"48",x"66",x"cc",x"87"),
  1481 => (x"a6",x"d0",x"88",x"c1"),
  1482 => (x"87",x"ce",x"c5",x"58"),
  1483 => (x"87",x"f6",x"d8",x"ff"),
  1484 => (x"58",x"a6",x"e8",x"c0"),
  1485 => (x"87",x"ee",x"d8",x"ff"),
  1486 => (x"58",x"a6",x"e0",x"c0"),
  1487 => (x"05",x"a8",x"ec",x"c0"),
  1488 => (x"dc",x"87",x"ca",x"c0"),
  1489 => (x"e4",x"c0",x"48",x"a6"),
  1490 => (x"c4",x"c0",x"78",x"66"),
  1491 => (x"e2",x"d5",x"ff",x"87"),
  1492 => (x"49",x"66",x"c8",x"87"),
  1493 => (x"fc",x"c0",x"91",x"cb"),
  1494 => (x"80",x"71",x"48",x"66"),
  1495 => (x"c8",x"4a",x"7e",x"70"),
  1496 => (x"ca",x"49",x"6e",x"82"),
  1497 => (x"66",x"e4",x"c0",x"81"),
  1498 => (x"49",x"66",x"dc",x"51"),
  1499 => (x"e4",x"c0",x"81",x"c1"),
  1500 => (x"48",x"c1",x"89",x"66"),
  1501 => (x"49",x"70",x"30",x"71"),
  1502 => (x"97",x"71",x"89",x"c1"),
  1503 => (x"c8",x"f9",x"c2",x"7a"),
  1504 => (x"e4",x"c0",x"49",x"bf"),
  1505 => (x"6a",x"97",x"29",x"66"),
  1506 => (x"98",x"71",x"48",x"4a"),
  1507 => (x"58",x"a6",x"ec",x"c0"),
  1508 => (x"81",x"c4",x"49",x"6e"),
  1509 => (x"66",x"d8",x"4d",x"69"),
  1510 => (x"a8",x"66",x"c4",x"48"),
  1511 => (x"87",x"c8",x"c0",x"02"),
  1512 => (x"c0",x"48",x"a6",x"c4"),
  1513 => (x"87",x"c5",x"c0",x"78"),
  1514 => (x"c1",x"48",x"a6",x"c4"),
  1515 => (x"1e",x"66",x"c4",x"78"),
  1516 => (x"75",x"1e",x"e0",x"c0"),
  1517 => (x"fe",x"d4",x"ff",x"49"),
  1518 => (x"70",x"86",x"c8",x"87"),
  1519 => (x"ac",x"b7",x"c0",x"4c"),
  1520 => (x"87",x"d4",x"c1",x"06"),
  1521 => (x"e0",x"c0",x"85",x"74"),
  1522 => (x"75",x"89",x"74",x"49"),
  1523 => (x"f5",x"e3",x"c1",x"4b"),
  1524 => (x"e3",x"fe",x"71",x"4a"),
  1525 => (x"85",x"c2",x"87",x"d1"),
  1526 => (x"48",x"66",x"e0",x"c0"),
  1527 => (x"e4",x"c0",x"80",x"c1"),
  1528 => (x"e8",x"c0",x"58",x"a6"),
  1529 => (x"81",x"c1",x"49",x"66"),
  1530 => (x"c0",x"02",x"a9",x"70"),
  1531 => (x"a6",x"c4",x"87",x"c8"),
  1532 => (x"c0",x"78",x"c0",x"48"),
  1533 => (x"a6",x"c4",x"87",x"c5"),
  1534 => (x"c4",x"78",x"c1",x"48"),
  1535 => (x"a4",x"c2",x"1e",x"66"),
  1536 => (x"48",x"e0",x"c0",x"49"),
  1537 => (x"49",x"70",x"88",x"71"),
  1538 => (x"ff",x"49",x"75",x"1e"),
  1539 => (x"c8",x"87",x"e8",x"d3"),
  1540 => (x"a8",x"b7",x"c0",x"86"),
  1541 => (x"87",x"c0",x"ff",x"01"),
  1542 => (x"02",x"66",x"e0",x"c0"),
  1543 => (x"6e",x"87",x"d1",x"c0"),
  1544 => (x"c0",x"81",x"c9",x"49"),
  1545 => (x"6e",x"51",x"66",x"e0"),
  1546 => (x"e3",x"cb",x"c1",x"48"),
  1547 => (x"87",x"cc",x"c0",x"78"),
  1548 => (x"81",x"c9",x"49",x"6e"),
  1549 => (x"48",x"6e",x"51",x"c2"),
  1550 => (x"78",x"cf",x"cd",x"c1"),
  1551 => (x"cc",x"48",x"66",x"c8"),
  1552 => (x"c0",x"04",x"a8",x"66"),
  1553 => (x"66",x"c8",x"87",x"cb"),
  1554 => (x"cc",x"80",x"c1",x"48"),
  1555 => (x"e9",x"c0",x"58",x"a6"),
  1556 => (x"48",x"66",x"cc",x"87"),
  1557 => (x"a6",x"d0",x"88",x"c1"),
  1558 => (x"87",x"de",x"c0",x"58"),
  1559 => (x"87",x"c3",x"d2",x"ff"),
  1560 => (x"d5",x"c0",x"4c",x"70"),
  1561 => (x"ac",x"c6",x"c1",x"87"),
  1562 => (x"87",x"c8",x"c0",x"05"),
  1563 => (x"c1",x"48",x"66",x"d0"),
  1564 => (x"58",x"a6",x"d4",x"80"),
  1565 => (x"87",x"eb",x"d1",x"ff"),
  1566 => (x"66",x"d4",x"4c",x"70"),
  1567 => (x"d8",x"80",x"c1",x"48"),
  1568 => (x"9c",x"74",x"58",x"a6"),
  1569 => (x"87",x"cb",x"c0",x"02"),
  1570 => (x"c1",x"48",x"66",x"c8"),
  1571 => (x"04",x"a8",x"66",x"c4"),
  1572 => (x"ff",x"87",x"f7",x"f2"),
  1573 => (x"c8",x"87",x"c3",x"d1"),
  1574 => (x"a8",x"c7",x"48",x"66"),
  1575 => (x"87",x"e5",x"c0",x"03"),
  1576 => (x"48",x"dc",x"f5",x"c2"),
  1577 => (x"66",x"c8",x"78",x"c0"),
  1578 => (x"c0",x"91",x"cb",x"49"),
  1579 => (x"c4",x"81",x"66",x"fc"),
  1580 => (x"4a",x"6a",x"4a",x"a1"),
  1581 => (x"c8",x"79",x"52",x"c0"),
  1582 => (x"80",x"c1",x"48",x"66"),
  1583 => (x"c7",x"58",x"a6",x"cc"),
  1584 => (x"db",x"ff",x"04",x"a8"),
  1585 => (x"8e",x"d4",x"ff",x"87"),
  1586 => (x"87",x"e9",x"db",x"ff"),
  1587 => (x"64",x"61",x"6f",x"4c"),
  1588 => (x"74",x"65",x"53",x"20"),
  1589 => (x"67",x"6e",x"69",x"74"),
  1590 => (x"00",x"81",x"20",x"73"),
  1591 => (x"65",x"76",x"61",x"53"),
  1592 => (x"74",x"65",x"53",x"20"),
  1593 => (x"67",x"6e",x"69",x"74"),
  1594 => (x"00",x"81",x"20",x"73"),
  1595 => (x"64",x"61",x"6f",x"4c"),
  1596 => (x"20",x"2e",x"2a",x"20"),
  1597 => (x"00",x"20",x"3a",x"00"),
  1598 => (x"71",x"1e",x"73",x"1e"),
  1599 => (x"c6",x"02",x"9b",x"4b"),
  1600 => (x"d8",x"f5",x"c2",x"87"),
  1601 => (x"c7",x"78",x"c0",x"48"),
  1602 => (x"d8",x"f5",x"c2",x"1e"),
  1603 => (x"e8",x"c1",x"1e",x"bf"),
  1604 => (x"f5",x"c2",x"1e",x"c3"),
  1605 => (x"eb",x"49",x"bf",x"c0"),
  1606 => (x"86",x"cc",x"87",x"e4"),
  1607 => (x"bf",x"c0",x"f5",x"c2"),
  1608 => (x"87",x"cd",x"e0",x"49"),
  1609 => (x"c8",x"02",x"9b",x"73"),
  1610 => (x"c3",x"e8",x"c1",x"87"),
  1611 => (x"c8",x"e2",x"c0",x"49"),
  1612 => (x"c4",x"da",x"ff",x"87"),
  1613 => (x"c1",x"c8",x"1e",x"87"),
  1614 => (x"fe",x"49",x"c1",x"87"),
  1615 => (x"f5",x"c2",x"87",x"fa"),
  1616 => (x"50",x"c0",x"48",x"e0"),
  1617 => (x"87",x"cf",x"e6",x"fe"),
  1618 => (x"cd",x"02",x"98",x"70"),
  1619 => (x"c9",x"ef",x"fe",x"87"),
  1620 => (x"02",x"98",x"70",x"87"),
  1621 => (x"4a",x"c1",x"87",x"c4"),
  1622 => (x"4a",x"c0",x"87",x"c2"),
  1623 => (x"ce",x"05",x"9a",x"72"),
  1624 => (x"c1",x"1e",x"c0",x"87"),
  1625 => (x"c0",x"49",x"ea",x"e6"),
  1626 => (x"c4",x"87",x"c5",x"f2"),
  1627 => (x"c1",x"87",x"fe",x"86"),
  1628 => (x"c0",x"49",x"f5",x"e6"),
  1629 => (x"c2",x"87",x"c7",x"fc"),
  1630 => (x"c0",x"48",x"d8",x"f5"),
  1631 => (x"c0",x"f5",x"c2",x"78"),
  1632 => (x"1e",x"78",x"c0",x"48"),
  1633 => (x"49",x"c1",x"e7",x"c1"),
  1634 => (x"87",x"e4",x"f1",x"c0"),
  1635 => (x"ff",x"c0",x"1e",x"c0"),
  1636 => (x"49",x"70",x"87",x"d1"),
  1637 => (x"87",x"d8",x"f1",x"c0"),
  1638 => (x"dc",x"c3",x"86",x"c8"),
  1639 => (x"db",x"e2",x"c0",x"87"),
  1640 => (x"da",x"f5",x"c0",x"87"),
  1641 => (x"87",x"f5",x"ff",x"87"),
  1642 => (x"44",x"53",x"4f",x"26"),
  1643 => (x"69",x"61",x"66",x"20"),
  1644 => (x"2e",x"64",x"65",x"6c"),
  1645 => (x"43",x"49",x"56",x"00"),
  1646 => (x"20",x"20",x"30",x"32"),
  1647 => (x"47",x"46",x"43",x"20"),
  1648 => (x"6f",x"6f",x"42",x"00"),
  1649 => (x"67",x"6e",x"69",x"74"),
  1650 => (x"00",x"2e",x"2e",x"2e"),
  1651 => (x"00",x"01",x"00",x"00"),
  1652 => (x"20",x"20",x"00",x"00"),
  1653 => (x"20",x"20",x"20",x"20"),
  1654 => (x"20",x"20",x"20",x"20"),
  1655 => (x"45",x"20",x"20",x"20"),
  1656 => (x"20",x"74",x"69",x"78"),
  1657 => (x"20",x"20",x"20",x"20"),
  1658 => (x"20",x"20",x"20",x"20"),
  1659 => (x"81",x"20",x"20",x"20"),
  1660 => (x"20",x"20",x"80",x"00"),
  1661 => (x"20",x"20",x"20",x"20"),
  1662 => (x"20",x"20",x"20",x"20"),
  1663 => (x"61",x"42",x"20",x"20"),
  1664 => (x"5e",x"00",x"6b",x"63"),
  1665 => (x"6c",x"00",x"00",x"10"),
  1666 => (x"00",x"00",x"00",x"2d"),
  1667 => (x"10",x"5e",x"00",x"00"),
  1668 => (x"2d",x"8a",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"00",x"10",x"5e",x"00"),
  1671 => (x"00",x"2d",x"a8",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"10",x"5e"),
  1674 => (x"00",x"00",x"2d",x"c6"),
  1675 => (x"5e",x"00",x"00",x"00"),
  1676 => (x"e4",x"00",x"00",x"10"),
  1677 => (x"00",x"00",x"00",x"2d"),
  1678 => (x"10",x"5e",x"00",x"00"),
  1679 => (x"2e",x"02",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"10",x"5e",x"00"),
  1682 => (x"00",x"2e",x"20",x"00"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"00",x"00",x"11",x"12"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"60",x"00",x"00",x"00"),
  1687 => (x"00",x"00",x"00",x"13"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"fe",x"1e",x"00",x"00"),
  1690 => (x"78",x"c0",x"48",x"f0"),
  1691 => (x"09",x"79",x"09",x"cd"),
  1692 => (x"fe",x"1e",x"4f",x"26"),
  1693 => (x"26",x"48",x"bf",x"f0"),
  1694 => (x"f0",x"fe",x"1e",x"4f"),
  1695 => (x"26",x"78",x"c1",x"48"),
  1696 => (x"f0",x"fe",x"1e",x"4f"),
  1697 => (x"26",x"78",x"c0",x"48"),
  1698 => (x"4a",x"71",x"1e",x"4f"),
  1699 => (x"26",x"51",x"52",x"c0"),
  1700 => (x"5b",x"5e",x"0e",x"4f"),
  1701 => (x"f4",x"0e",x"5d",x"5c"),
  1702 => (x"97",x"4d",x"71",x"86"),
  1703 => (x"a5",x"c1",x"7e",x"6d"),
  1704 => (x"48",x"6c",x"97",x"4c"),
  1705 => (x"6e",x"58",x"a6",x"c8"),
  1706 => (x"a8",x"66",x"c4",x"48"),
  1707 => (x"ff",x"87",x"c5",x"05"),
  1708 => (x"87",x"e6",x"c0",x"48"),
  1709 => (x"c2",x"87",x"ca",x"ff"),
  1710 => (x"6c",x"97",x"49",x"a5"),
  1711 => (x"4b",x"a3",x"71",x"4b"),
  1712 => (x"97",x"4b",x"6b",x"97"),
  1713 => (x"48",x"6e",x"7e",x"6c"),
  1714 => (x"a6",x"c8",x"80",x"c1"),
  1715 => (x"cc",x"98",x"c7",x"58"),
  1716 => (x"97",x"70",x"58",x"a6"),
  1717 => (x"87",x"e1",x"fe",x"7c"),
  1718 => (x"8e",x"f4",x"48",x"73"),
  1719 => (x"4c",x"26",x"4d",x"26"),
  1720 => (x"4f",x"26",x"4b",x"26"),
  1721 => (x"5c",x"5b",x"5e",x"0e"),
  1722 => (x"71",x"86",x"f4",x"0e"),
  1723 => (x"4a",x"66",x"d8",x"4c"),
  1724 => (x"c2",x"9a",x"ff",x"c3"),
  1725 => (x"6c",x"97",x"4b",x"a4"),
  1726 => (x"49",x"a1",x"73",x"49"),
  1727 => (x"6c",x"97",x"51",x"72"),
  1728 => (x"c1",x"48",x"6e",x"7e"),
  1729 => (x"58",x"a6",x"c8",x"80"),
  1730 => (x"a6",x"cc",x"98",x"c7"),
  1731 => (x"f4",x"54",x"70",x"58"),
  1732 => (x"87",x"ca",x"ff",x"8e"),
  1733 => (x"e8",x"fd",x"1e",x"1e"),
  1734 => (x"4a",x"bf",x"e0",x"87"),
  1735 => (x"c0",x"e0",x"c0",x"49"),
  1736 => (x"87",x"cb",x"02",x"99"),
  1737 => (x"f8",x"c2",x"1e",x"72"),
  1738 => (x"f7",x"fe",x"49",x"fe"),
  1739 => (x"fd",x"86",x"c4",x"87"),
  1740 => (x"7e",x"70",x"87",x"c0"),
  1741 => (x"26",x"87",x"c2",x"fd"),
  1742 => (x"c2",x"1e",x"4f",x"26"),
  1743 => (x"fd",x"49",x"fe",x"f8"),
  1744 => (x"ec",x"c1",x"87",x"c7"),
  1745 => (x"dd",x"fc",x"49",x"d4"),
  1746 => (x"87",x"f5",x"c2",x"87"),
  1747 => (x"73",x"1e",x"4f",x"26"),
  1748 => (x"fe",x"f8",x"c2",x"1e"),
  1749 => (x"87",x"f9",x"fc",x"49"),
  1750 => (x"b7",x"c0",x"4a",x"70"),
  1751 => (x"cc",x"c2",x"04",x"aa"),
  1752 => (x"aa",x"f0",x"c3",x"87"),
  1753 => (x"c1",x"87",x"c9",x"05"),
  1754 => (x"c1",x"48",x"f9",x"ef"),
  1755 => (x"87",x"ed",x"c1",x"78"),
  1756 => (x"05",x"aa",x"e0",x"c3"),
  1757 => (x"ef",x"c1",x"87",x"c9"),
  1758 => (x"78",x"c1",x"48",x"fd"),
  1759 => (x"c1",x"87",x"de",x"c1"),
  1760 => (x"02",x"bf",x"fd",x"ef"),
  1761 => (x"c0",x"c2",x"87",x"c6"),
  1762 => (x"87",x"c2",x"4b",x"a2"),
  1763 => (x"ef",x"c1",x"4b",x"72"),
  1764 => (x"c0",x"02",x"bf",x"f9"),
  1765 => (x"49",x"73",x"87",x"e0"),
  1766 => (x"91",x"29",x"b7",x"c4"),
  1767 => (x"81",x"d0",x"f1",x"c1"),
  1768 => (x"9a",x"cf",x"4a",x"73"),
  1769 => (x"48",x"c1",x"92",x"c2"),
  1770 => (x"4a",x"70",x"30",x"72"),
  1771 => (x"48",x"72",x"ba",x"ff"),
  1772 => (x"79",x"70",x"98",x"69"),
  1773 => (x"49",x"73",x"87",x"db"),
  1774 => (x"91",x"29",x"b7",x"c4"),
  1775 => (x"81",x"d0",x"f1",x"c1"),
  1776 => (x"9a",x"cf",x"4a",x"73"),
  1777 => (x"48",x"c3",x"92",x"c2"),
  1778 => (x"4a",x"70",x"30",x"72"),
  1779 => (x"70",x"b0",x"69",x"48"),
  1780 => (x"fd",x"ef",x"c1",x"79"),
  1781 => (x"c1",x"78",x"c0",x"48"),
  1782 => (x"c0",x"48",x"f9",x"ef"),
  1783 => (x"fe",x"f8",x"c2",x"78"),
  1784 => (x"87",x"ed",x"fa",x"49"),
  1785 => (x"b7",x"c0",x"4a",x"70"),
  1786 => (x"f4",x"fd",x"03",x"aa"),
  1787 => (x"c4",x"48",x"c0",x"87"),
  1788 => (x"26",x"4d",x"26",x"87"),
  1789 => (x"26",x"4b",x"26",x"4c"),
  1790 => (x"00",x"00",x"00",x"4f"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"4a",x"c0",x"1e",x"00"),
  1793 => (x"91",x"c4",x"49",x"72"),
  1794 => (x"81",x"d0",x"f1",x"c1"),
  1795 => (x"82",x"c1",x"79",x"c0"),
  1796 => (x"04",x"aa",x"b7",x"d0"),
  1797 => (x"4f",x"26",x"87",x"ee"),
  1798 => (x"5c",x"5b",x"5e",x"0e"),
  1799 => (x"4d",x"71",x"0e",x"5d"),
  1800 => (x"75",x"87",x"de",x"f9"),
  1801 => (x"2a",x"b7",x"c4",x"4a"),
  1802 => (x"d0",x"f1",x"c1",x"92"),
  1803 => (x"cf",x"4c",x"75",x"82"),
  1804 => (x"6a",x"94",x"c2",x"9c"),
  1805 => (x"2b",x"74",x"4b",x"49"),
  1806 => (x"48",x"c2",x"9b",x"c3"),
  1807 => (x"4c",x"70",x"30",x"74"),
  1808 => (x"48",x"74",x"bc",x"ff"),
  1809 => (x"7a",x"70",x"98",x"71"),
  1810 => (x"73",x"87",x"ee",x"f8"),
  1811 => (x"87",x"e1",x"fe",x"48"),
  1812 => (x"00",x"00",x"00",x"00"),
  1813 => (x"00",x"00",x"00",x"00"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"00",x"00",x"00",x"00"),
  1816 => (x"00",x"00",x"00",x"00"),
  1817 => (x"00",x"00",x"00",x"00"),
  1818 => (x"00",x"00",x"00",x"00"),
  1819 => (x"00",x"00",x"00",x"00"),
  1820 => (x"00",x"00",x"00",x"00"),
  1821 => (x"00",x"00",x"00",x"00"),
  1822 => (x"00",x"00",x"00",x"00"),
  1823 => (x"00",x"00",x"00",x"00"),
  1824 => (x"00",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"48",x"d0",x"ff",x"1e"),
  1829 => (x"71",x"78",x"e1",x"c8"),
  1830 => (x"08",x"d4",x"ff",x"48"),
  1831 => (x"1e",x"4f",x"26",x"78"),
  1832 => (x"c8",x"48",x"d0",x"ff"),
  1833 => (x"48",x"71",x"78",x"e1"),
  1834 => (x"78",x"08",x"d4",x"ff"),
  1835 => (x"ff",x"48",x"66",x"c4"),
  1836 => (x"26",x"78",x"08",x"d4"),
  1837 => (x"4a",x"71",x"1e",x"4f"),
  1838 => (x"1e",x"49",x"66",x"c4"),
  1839 => (x"de",x"ff",x"49",x"72"),
  1840 => (x"48",x"d0",x"ff",x"87"),
  1841 => (x"26",x"78",x"e0",x"c0"),
  1842 => (x"73",x"1e",x"4f",x"26"),
  1843 => (x"c8",x"4b",x"71",x"1e"),
  1844 => (x"73",x"1e",x"49",x"66"),
  1845 => (x"a2",x"e0",x"c1",x"4a"),
  1846 => (x"87",x"d9",x"ff",x"49"),
  1847 => (x"26",x"87",x"c4",x"26"),
  1848 => (x"26",x"4c",x"26",x"4d"),
  1849 => (x"1e",x"4f",x"26",x"4b"),
  1850 => (x"c3",x"4a",x"d4",x"ff"),
  1851 => (x"d0",x"ff",x"7a",x"ff"),
  1852 => (x"78",x"e1",x"c0",x"48"),
  1853 => (x"f9",x"c2",x"7a",x"de"),
  1854 => (x"49",x"7a",x"bf",x"c8"),
  1855 => (x"70",x"28",x"c8",x"48"),
  1856 => (x"d0",x"48",x"71",x"7a"),
  1857 => (x"71",x"7a",x"70",x"28"),
  1858 => (x"70",x"28",x"d8",x"48"),
  1859 => (x"48",x"d0",x"ff",x"7a"),
  1860 => (x"26",x"78",x"e0",x"c0"),
  1861 => (x"d0",x"ff",x"1e",x"4f"),
  1862 => (x"78",x"c9",x"c8",x"48"),
  1863 => (x"d4",x"ff",x"48",x"71"),
  1864 => (x"4f",x"26",x"78",x"08"),
  1865 => (x"49",x"4a",x"71",x"1e"),
  1866 => (x"d0",x"ff",x"87",x"eb"),
  1867 => (x"26",x"78",x"c8",x"48"),
  1868 => (x"1e",x"73",x"1e",x"4f"),
  1869 => (x"f9",x"c2",x"4b",x"71"),
  1870 => (x"c3",x"02",x"bf",x"d8"),
  1871 => (x"87",x"eb",x"c2",x"87"),
  1872 => (x"c8",x"48",x"d0",x"ff"),
  1873 => (x"48",x"73",x"78",x"c9"),
  1874 => (x"ff",x"b0",x"e0",x"c0"),
  1875 => (x"c2",x"78",x"08",x"d4"),
  1876 => (x"c0",x"48",x"cc",x"f9"),
  1877 => (x"02",x"66",x"c8",x"78"),
  1878 => (x"ff",x"c3",x"87",x"c5"),
  1879 => (x"c0",x"87",x"c2",x"49"),
  1880 => (x"d4",x"f9",x"c2",x"49"),
  1881 => (x"02",x"66",x"cc",x"59"),
  1882 => (x"d5",x"c5",x"87",x"c6"),
  1883 => (x"87",x"c4",x"4a",x"d5"),
  1884 => (x"4a",x"ff",x"ff",x"cf"),
  1885 => (x"5a",x"d8",x"f9",x"c2"),
  1886 => (x"48",x"d8",x"f9",x"c2"),
  1887 => (x"87",x"c4",x"78",x"c1"),
  1888 => (x"4c",x"26",x"4d",x"26"),
  1889 => (x"4f",x"26",x"4b",x"26"),
  1890 => (x"5c",x"5b",x"5e",x"0e"),
  1891 => (x"4a",x"71",x"0e",x"5d"),
  1892 => (x"bf",x"d4",x"f9",x"c2"),
  1893 => (x"02",x"9a",x"72",x"4c"),
  1894 => (x"c8",x"49",x"87",x"cb"),
  1895 => (x"e7",x"f4",x"c1",x"91"),
  1896 => (x"c4",x"83",x"71",x"4b"),
  1897 => (x"e7",x"f8",x"c1",x"87"),
  1898 => (x"13",x"4d",x"c0",x"4b"),
  1899 => (x"c2",x"99",x"74",x"49"),
  1900 => (x"48",x"bf",x"d0",x"f9"),
  1901 => (x"d4",x"ff",x"b8",x"71"),
  1902 => (x"b7",x"c1",x"78",x"08"),
  1903 => (x"b7",x"c8",x"85",x"2c"),
  1904 => (x"87",x"e7",x"04",x"ad"),
  1905 => (x"bf",x"cc",x"f9",x"c2"),
  1906 => (x"c2",x"80",x"c8",x"48"),
  1907 => (x"fe",x"58",x"d0",x"f9"),
  1908 => (x"73",x"1e",x"87",x"ee"),
  1909 => (x"13",x"4b",x"71",x"1e"),
  1910 => (x"cb",x"02",x"9a",x"4a"),
  1911 => (x"fe",x"49",x"72",x"87"),
  1912 => (x"4a",x"13",x"87",x"e6"),
  1913 => (x"87",x"f5",x"05",x"9a"),
  1914 => (x"1e",x"87",x"d9",x"fe"),
  1915 => (x"bf",x"cc",x"f9",x"c2"),
  1916 => (x"cc",x"f9",x"c2",x"49"),
  1917 => (x"78",x"a1",x"c1",x"48"),
  1918 => (x"a9",x"b7",x"c0",x"c4"),
  1919 => (x"ff",x"87",x"db",x"03"),
  1920 => (x"f9",x"c2",x"48",x"d4"),
  1921 => (x"c2",x"78",x"bf",x"d0"),
  1922 => (x"49",x"bf",x"cc",x"f9"),
  1923 => (x"48",x"cc",x"f9",x"c2"),
  1924 => (x"c4",x"78",x"a1",x"c1"),
  1925 => (x"04",x"a9",x"b7",x"c0"),
  1926 => (x"d0",x"ff",x"87",x"e5"),
  1927 => (x"c2",x"78",x"c8",x"48"),
  1928 => (x"c0",x"48",x"d8",x"f9"),
  1929 => (x"00",x"4f",x"26",x"78"),
  1930 => (x"00",x"00",x"00",x"00"),
  1931 => (x"00",x"00",x"00",x"00"),
  1932 => (x"5f",x"5f",x"00",x"00"),
  1933 => (x"00",x"00",x"00",x"00"),
  1934 => (x"03",x"00",x"03",x"03"),
  1935 => (x"14",x"00",x"00",x"03"),
  1936 => (x"7f",x"14",x"7f",x"7f"),
  1937 => (x"00",x"00",x"14",x"7f"),
  1938 => (x"6b",x"6b",x"2e",x"24"),
  1939 => (x"4c",x"00",x"12",x"3a"),
  1940 => (x"6c",x"18",x"36",x"6a"),
  1941 => (x"30",x"00",x"32",x"56"),
  1942 => (x"77",x"59",x"4f",x"7e"),
  1943 => (x"00",x"40",x"68",x"3a"),
  1944 => (x"03",x"07",x"04",x"00"),
  1945 => (x"00",x"00",x"00",x"00"),
  1946 => (x"63",x"3e",x"1c",x"00"),
  1947 => (x"00",x"00",x"00",x"41"),
  1948 => (x"3e",x"63",x"41",x"00"),
  1949 => (x"08",x"00",x"00",x"1c"),
  1950 => (x"1c",x"1c",x"3e",x"2a"),
  1951 => (x"00",x"08",x"2a",x"3e"),
  1952 => (x"3e",x"3e",x"08",x"08"),
  1953 => (x"00",x"00",x"08",x"08"),
  1954 => (x"60",x"e0",x"80",x"00"),
  1955 => (x"00",x"00",x"00",x"00"),
  1956 => (x"08",x"08",x"08",x"08"),
  1957 => (x"00",x"00",x"08",x"08"),
  1958 => (x"60",x"60",x"00",x"00"),
  1959 => (x"40",x"00",x"00",x"00"),
  1960 => (x"0c",x"18",x"30",x"60"),
  1961 => (x"00",x"01",x"03",x"06"),
  1962 => (x"4d",x"59",x"7f",x"3e"),
  1963 => (x"00",x"00",x"3e",x"7f"),
  1964 => (x"7f",x"7f",x"06",x"04"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"59",x"71",x"63",x"42"),
  1967 => (x"00",x"00",x"46",x"4f"),
  1968 => (x"49",x"49",x"63",x"22"),
  1969 => (x"18",x"00",x"36",x"7f"),
  1970 => (x"7f",x"13",x"16",x"1c"),
  1971 => (x"00",x"00",x"10",x"7f"),
  1972 => (x"45",x"45",x"67",x"27"),
  1973 => (x"00",x"00",x"39",x"7d"),
  1974 => (x"49",x"4b",x"7e",x"3c"),
  1975 => (x"00",x"00",x"30",x"79"),
  1976 => (x"79",x"71",x"01",x"01"),
  1977 => (x"00",x"00",x"07",x"0f"),
  1978 => (x"49",x"49",x"7f",x"36"),
  1979 => (x"00",x"00",x"36",x"7f"),
  1980 => (x"69",x"49",x"4f",x"06"),
  1981 => (x"00",x"00",x"1e",x"3f"),
  1982 => (x"66",x"66",x"00",x"00"),
  1983 => (x"00",x"00",x"00",x"00"),
  1984 => (x"66",x"e6",x"80",x"00"),
  1985 => (x"00",x"00",x"00",x"00"),
  1986 => (x"14",x"14",x"08",x"08"),
  1987 => (x"00",x"00",x"22",x"22"),
  1988 => (x"14",x"14",x"14",x"14"),
  1989 => (x"00",x"00",x"14",x"14"),
  1990 => (x"14",x"14",x"22",x"22"),
  1991 => (x"00",x"00",x"08",x"08"),
  1992 => (x"59",x"51",x"03",x"02"),
  1993 => (x"3e",x"00",x"06",x"0f"),
  1994 => (x"55",x"5d",x"41",x"7f"),
  1995 => (x"00",x"00",x"1e",x"1f"),
  1996 => (x"09",x"09",x"7f",x"7e"),
  1997 => (x"00",x"00",x"7e",x"7f"),
  1998 => (x"49",x"49",x"7f",x"7f"),
  1999 => (x"00",x"00",x"36",x"7f"),
  2000 => (x"41",x"63",x"3e",x"1c"),
  2001 => (x"00",x"00",x"41",x"41"),
  2002 => (x"63",x"41",x"7f",x"7f"),
  2003 => (x"00",x"00",x"1c",x"3e"),
  2004 => (x"49",x"49",x"7f",x"7f"),
  2005 => (x"00",x"00",x"41",x"41"),
  2006 => (x"09",x"09",x"7f",x"7f"),
  2007 => (x"00",x"00",x"01",x"01"),
  2008 => (x"49",x"41",x"7f",x"3e"),
  2009 => (x"00",x"00",x"7a",x"7b"),
  2010 => (x"08",x"08",x"7f",x"7f"),
  2011 => (x"00",x"00",x"7f",x"7f"),
  2012 => (x"7f",x"7f",x"41",x"00"),
  2013 => (x"00",x"00",x"00",x"41"),
  2014 => (x"40",x"40",x"60",x"20"),
  2015 => (x"7f",x"00",x"3f",x"7f"),
  2016 => (x"36",x"1c",x"08",x"7f"),
  2017 => (x"00",x"00",x"41",x"63"),
  2018 => (x"40",x"40",x"7f",x"7f"),
  2019 => (x"7f",x"00",x"40",x"40"),
  2020 => (x"06",x"0c",x"06",x"7f"),
  2021 => (x"7f",x"00",x"7f",x"7f"),
  2022 => (x"18",x"0c",x"06",x"7f"),
  2023 => (x"00",x"00",x"7f",x"7f"),
  2024 => (x"41",x"41",x"7f",x"3e"),
  2025 => (x"00",x"00",x"3e",x"7f"),
  2026 => (x"09",x"09",x"7f",x"7f"),
  2027 => (x"3e",x"00",x"06",x"0f"),
  2028 => (x"7f",x"61",x"41",x"7f"),
  2029 => (x"00",x"00",x"40",x"7e"),
  2030 => (x"19",x"09",x"7f",x"7f"),
  2031 => (x"00",x"00",x"66",x"7f"),
  2032 => (x"59",x"4d",x"6f",x"26"),
  2033 => (x"00",x"00",x"32",x"7b"),
  2034 => (x"7f",x"7f",x"01",x"01"),
  2035 => (x"00",x"00",x"01",x"01"),
  2036 => (x"40",x"40",x"7f",x"3f"),
  2037 => (x"00",x"00",x"3f",x"7f"),
  2038 => (x"70",x"70",x"3f",x"0f"),
  2039 => (x"7f",x"00",x"0f",x"3f"),
  2040 => (x"30",x"18",x"30",x"7f"),
  2041 => (x"41",x"00",x"7f",x"7f"),
  2042 => (x"1c",x"1c",x"36",x"63"),
  2043 => (x"01",x"41",x"63",x"36"),
  2044 => (x"7c",x"7c",x"06",x"03"),
  2045 => (x"61",x"01",x"03",x"06"),
  2046 => (x"47",x"4d",x"59",x"71"),
  2047 => (x"00",x"00",x"41",x"43"),
  2048 => (x"41",x"7f",x"7f",x"00"),
  2049 => (x"01",x"00",x"00",x"41"),
  2050 => (x"18",x"0c",x"06",x"03"),
  2051 => (x"00",x"40",x"60",x"30"),
  2052 => (x"7f",x"41",x"41",x"00"),
  2053 => (x"08",x"00",x"00",x"7f"),
  2054 => (x"06",x"03",x"06",x"0c"),
  2055 => (x"80",x"00",x"08",x"0c"),
  2056 => (x"80",x"80",x"80",x"80"),
  2057 => (x"00",x"00",x"80",x"80"),
  2058 => (x"07",x"03",x"00",x"00"),
  2059 => (x"00",x"00",x"00",x"04"),
  2060 => (x"54",x"54",x"74",x"20"),
  2061 => (x"00",x"00",x"78",x"7c"),
  2062 => (x"44",x"44",x"7f",x"7f"),
  2063 => (x"00",x"00",x"38",x"7c"),
  2064 => (x"44",x"44",x"7c",x"38"),
  2065 => (x"00",x"00",x"00",x"44"),
  2066 => (x"44",x"44",x"7c",x"38"),
  2067 => (x"00",x"00",x"7f",x"7f"),
  2068 => (x"54",x"54",x"7c",x"38"),
  2069 => (x"00",x"00",x"18",x"5c"),
  2070 => (x"05",x"7f",x"7e",x"04"),
  2071 => (x"00",x"00",x"00",x"05"),
  2072 => (x"a4",x"a4",x"bc",x"18"),
  2073 => (x"00",x"00",x"7c",x"fc"),
  2074 => (x"04",x"04",x"7f",x"7f"),
  2075 => (x"00",x"00",x"78",x"7c"),
  2076 => (x"7d",x"3d",x"00",x"00"),
  2077 => (x"00",x"00",x"00",x"40"),
  2078 => (x"fd",x"80",x"80",x"80"),
  2079 => (x"00",x"00",x"00",x"7d"),
  2080 => (x"38",x"10",x"7f",x"7f"),
  2081 => (x"00",x"00",x"44",x"6c"),
  2082 => (x"7f",x"3f",x"00",x"00"),
  2083 => (x"7c",x"00",x"00",x"40"),
  2084 => (x"0c",x"18",x"0c",x"7c"),
  2085 => (x"00",x"00",x"78",x"7c"),
  2086 => (x"04",x"04",x"7c",x"7c"),
  2087 => (x"00",x"00",x"78",x"7c"),
  2088 => (x"44",x"44",x"7c",x"38"),
  2089 => (x"00",x"00",x"38",x"7c"),
  2090 => (x"24",x"24",x"fc",x"fc"),
  2091 => (x"00",x"00",x"18",x"3c"),
  2092 => (x"24",x"24",x"3c",x"18"),
  2093 => (x"00",x"00",x"fc",x"fc"),
  2094 => (x"04",x"04",x"7c",x"7c"),
  2095 => (x"00",x"00",x"08",x"0c"),
  2096 => (x"54",x"54",x"5c",x"48"),
  2097 => (x"00",x"00",x"20",x"74"),
  2098 => (x"44",x"7f",x"3f",x"04"),
  2099 => (x"00",x"00",x"00",x"44"),
  2100 => (x"40",x"40",x"7c",x"3c"),
  2101 => (x"00",x"00",x"7c",x"7c"),
  2102 => (x"60",x"60",x"3c",x"1c"),
  2103 => (x"3c",x"00",x"1c",x"3c"),
  2104 => (x"60",x"30",x"60",x"7c"),
  2105 => (x"44",x"00",x"3c",x"7c"),
  2106 => (x"38",x"10",x"38",x"6c"),
  2107 => (x"00",x"00",x"44",x"6c"),
  2108 => (x"60",x"e0",x"bc",x"1c"),
  2109 => (x"00",x"00",x"1c",x"3c"),
  2110 => (x"5c",x"74",x"64",x"44"),
  2111 => (x"00",x"00",x"44",x"4c"),
  2112 => (x"77",x"3e",x"08",x"08"),
  2113 => (x"00",x"00",x"41",x"41"),
  2114 => (x"7f",x"7f",x"00",x"00"),
  2115 => (x"00",x"00",x"00",x"00"),
  2116 => (x"3e",x"77",x"41",x"41"),
  2117 => (x"02",x"00",x"08",x"08"),
  2118 => (x"02",x"03",x"01",x"01"),
  2119 => (x"7f",x"00",x"01",x"02"),
  2120 => (x"7f",x"7f",x"7f",x"7f"),
  2121 => (x"08",x"00",x"7f",x"7f"),
  2122 => (x"3e",x"1c",x"1c",x"08"),
  2123 => (x"7f",x"7f",x"7f",x"3e"),
  2124 => (x"1c",x"3e",x"3e",x"7f"),
  2125 => (x"00",x"08",x"08",x"1c"),
  2126 => (x"7c",x"7c",x"18",x"10"),
  2127 => (x"00",x"00",x"10",x"18"),
  2128 => (x"7c",x"7c",x"30",x"10"),
  2129 => (x"10",x"00",x"10",x"30"),
  2130 => (x"78",x"60",x"60",x"30"),
  2131 => (x"42",x"00",x"06",x"1e"),
  2132 => (x"3c",x"18",x"3c",x"66"),
  2133 => (x"78",x"00",x"42",x"66"),
  2134 => (x"c6",x"c2",x"6a",x"38"),
  2135 => (x"60",x"00",x"38",x"6c"),
  2136 => (x"00",x"60",x"00",x"00"),
  2137 => (x"0e",x"00",x"60",x"00"),
  2138 => (x"5d",x"5c",x"5b",x"5e"),
  2139 => (x"4c",x"71",x"1e",x"0e"),
  2140 => (x"bf",x"dd",x"f9",x"c2"),
  2141 => (x"c0",x"4b",x"c0",x"4d"),
  2142 => (x"02",x"ab",x"74",x"1e"),
  2143 => (x"a6",x"c4",x"87",x"c7"),
  2144 => (x"c5",x"78",x"c0",x"48"),
  2145 => (x"48",x"a6",x"c4",x"87"),
  2146 => (x"66",x"c4",x"78",x"c1"),
  2147 => (x"ee",x"49",x"73",x"1e"),
  2148 => (x"86",x"c8",x"87",x"df"),
  2149 => (x"ef",x"49",x"e0",x"c0"),
  2150 => (x"a5",x"c4",x"87",x"ee"),
  2151 => (x"f0",x"49",x"6a",x"4a"),
  2152 => (x"c6",x"f1",x"87",x"f0"),
  2153 => (x"c1",x"85",x"cb",x"87"),
  2154 => (x"ab",x"b7",x"c8",x"83"),
  2155 => (x"87",x"c7",x"ff",x"04"),
  2156 => (x"26",x"4d",x"26",x"26"),
  2157 => (x"26",x"4b",x"26",x"4c"),
  2158 => (x"4a",x"71",x"1e",x"4f"),
  2159 => (x"5a",x"e1",x"f9",x"c2"),
  2160 => (x"48",x"e1",x"f9",x"c2"),
  2161 => (x"fe",x"49",x"78",x"c7"),
  2162 => (x"4f",x"26",x"87",x"dd"),
  2163 => (x"71",x"1e",x"73",x"1e"),
  2164 => (x"aa",x"b7",x"c0",x"4a"),
  2165 => (x"c2",x"87",x"d3",x"03"),
  2166 => (x"05",x"bf",x"de",x"d9"),
  2167 => (x"4b",x"c1",x"87",x"c4"),
  2168 => (x"4b",x"c0",x"87",x"c2"),
  2169 => (x"5b",x"e2",x"d9",x"c2"),
  2170 => (x"d9",x"c2",x"87",x"c4"),
  2171 => (x"d9",x"c2",x"5a",x"e2"),
  2172 => (x"c1",x"4a",x"bf",x"de"),
  2173 => (x"a2",x"c0",x"c1",x"9a"),
  2174 => (x"87",x"e8",x"ec",x"49"),
  2175 => (x"bf",x"c6",x"d9",x"c2"),
  2176 => (x"de",x"d9",x"c2",x"48"),
  2177 => (x"08",x"fc",x"b0",x"bf"),
  2178 => (x"87",x"e9",x"fe",x"78"),
  2179 => (x"c4",x"4a",x"71",x"1e"),
  2180 => (x"49",x"72",x"1e",x"66"),
  2181 => (x"26",x"87",x"f3",x"ea"),
  2182 => (x"ff",x"1e",x"4f",x"26"),
  2183 => (x"ff",x"c3",x"48",x"d4"),
  2184 => (x"48",x"d0",x"ff",x"78"),
  2185 => (x"ff",x"78",x"e1",x"c0"),
  2186 => (x"78",x"c1",x"48",x"d4"),
  2187 => (x"30",x"c4",x"48",x"71"),
  2188 => (x"78",x"08",x"d4",x"ff"),
  2189 => (x"c0",x"48",x"d0",x"ff"),
  2190 => (x"4f",x"26",x"78",x"e0"),
  2191 => (x"5c",x"5b",x"5e",x"0e"),
  2192 => (x"86",x"f4",x"0e",x"5d"),
  2193 => (x"c0",x"48",x"a6",x"c4"),
  2194 => (x"bf",x"ec",x"4b",x"78"),
  2195 => (x"dd",x"f9",x"c2",x"7e"),
  2196 => (x"bf",x"e8",x"4d",x"bf"),
  2197 => (x"de",x"d9",x"c2",x"4c"),
  2198 => (x"f1",x"e3",x"49",x"bf"),
  2199 => (x"49",x"f7",x"c1",x"87"),
  2200 => (x"70",x"87",x"f5",x"e6"),
  2201 => (x"87",x"d5",x"02",x"98"),
  2202 => (x"bf",x"de",x"d9",x"c2"),
  2203 => (x"87",x"de",x"e3",x"49"),
  2204 => (x"f7",x"c1",x"4b",x"c1"),
  2205 => (x"87",x"e0",x"e6",x"49"),
  2206 => (x"eb",x"05",x"98",x"70"),
  2207 => (x"02",x"9b",x"73",x"87"),
  2208 => (x"c2",x"87",x"fa",x"c0"),
  2209 => (x"05",x"bf",x"c6",x"d9"),
  2210 => (x"a6",x"c8",x"87",x"c7"),
  2211 => (x"c5",x"78",x"c1",x"48"),
  2212 => (x"48",x"a6",x"c8",x"87"),
  2213 => (x"d9",x"c2",x"78",x"c0"),
  2214 => (x"66",x"c8",x"48",x"c6"),
  2215 => (x"1e",x"fc",x"ca",x"78"),
  2216 => (x"c9",x"02",x"66",x"cc"),
  2217 => (x"48",x"a6",x"cc",x"87"),
  2218 => (x"78",x"d9",x"d7",x"c2"),
  2219 => (x"a6",x"cc",x"87",x"c7"),
  2220 => (x"e4",x"d7",x"c2",x"48"),
  2221 => (x"49",x"66",x"cc",x"78"),
  2222 => (x"c4",x"87",x"f5",x"cc"),
  2223 => (x"cb",x"4b",x"c0",x"86"),
  2224 => (x"e1",x"ce",x"49",x"ee"),
  2225 => (x"58",x"a6",x"cc",x"87"),
  2226 => (x"cb",x"e5",x"49",x"c7"),
  2227 => (x"05",x"98",x"70",x"87"),
  2228 => (x"49",x"6e",x"87",x"c8"),
  2229 => (x"c1",x"02",x"99",x"c1"),
  2230 => (x"4b",x"c1",x"87",x"c3"),
  2231 => (x"c2",x"7e",x"bf",x"ec"),
  2232 => (x"49",x"bf",x"de",x"d9"),
  2233 => (x"c8",x"87",x"e7",x"e1"),
  2234 => (x"c5",x"ce",x"49",x"66"),
  2235 => (x"02",x"98",x"70",x"87"),
  2236 => (x"d9",x"c2",x"87",x"d8"),
  2237 => (x"c1",x"49",x"bf",x"c2"),
  2238 => (x"c6",x"d9",x"c2",x"b9"),
  2239 => (x"d9",x"fc",x"71",x"59"),
  2240 => (x"49",x"ee",x"cb",x"87"),
  2241 => (x"cc",x"87",x"df",x"cd"),
  2242 => (x"49",x"c7",x"58",x"a6"),
  2243 => (x"70",x"87",x"c9",x"e4"),
  2244 => (x"c5",x"ff",x"05",x"98"),
  2245 => (x"c1",x"49",x"6e",x"87"),
  2246 => (x"fd",x"fe",x"05",x"99"),
  2247 => (x"02",x"9b",x"73",x"87"),
  2248 => (x"49",x"ff",x"87",x"d0"),
  2249 => (x"c1",x"87",x"e5",x"fa"),
  2250 => (x"eb",x"e3",x"49",x"da"),
  2251 => (x"48",x"a6",x"c4",x"87"),
  2252 => (x"d9",x"c2",x"78",x"c1"),
  2253 => (x"c1",x"05",x"bf",x"de"),
  2254 => (x"d9",x"c2",x"87",x"e2"),
  2255 => (x"c0",x"02",x"bf",x"c6"),
  2256 => (x"a6",x"c4",x"87",x"f1"),
  2257 => (x"c0",x"c0",x"c8",x"48"),
  2258 => (x"ca",x"d9",x"c2",x"78"),
  2259 => (x"bf",x"97",x"6e",x"7e"),
  2260 => (x"c1",x"48",x"6e",x"49"),
  2261 => (x"71",x"7e",x"70",x"80"),
  2262 => (x"70",x"87",x"fd",x"e2"),
  2263 => (x"c3",x"c0",x"02",x"98"),
  2264 => (x"b4",x"66",x"c4",x"87"),
  2265 => (x"c1",x"48",x"66",x"c4"),
  2266 => (x"a6",x"c8",x"28",x"b7"),
  2267 => (x"05",x"98",x"70",x"58"),
  2268 => (x"c3",x"87",x"da",x"ff"),
  2269 => (x"df",x"e2",x"49",x"fd"),
  2270 => (x"49",x"fa",x"c3",x"87"),
  2271 => (x"74",x"87",x"d9",x"e2"),
  2272 => (x"99",x"ff",x"c3",x"49"),
  2273 => (x"49",x"c0",x"1e",x"71"),
  2274 => (x"74",x"87",x"c1",x"fa"),
  2275 => (x"29",x"b7",x"c8",x"49"),
  2276 => (x"49",x"c1",x"1e",x"71"),
  2277 => (x"c8",x"87",x"f5",x"f9"),
  2278 => (x"87",x"f8",x"c8",x"86"),
  2279 => (x"ff",x"c3",x"49",x"74"),
  2280 => (x"2c",x"b7",x"c8",x"99"),
  2281 => (x"9c",x"74",x"b4",x"71"),
  2282 => (x"87",x"e0",x"c0",x"02"),
  2283 => (x"bf",x"da",x"d9",x"c2"),
  2284 => (x"87",x"fe",x"ca",x"49"),
  2285 => (x"c0",x"05",x"98",x"70"),
  2286 => (x"4c",x"c0",x"87",x"c5"),
  2287 => (x"c2",x"87",x"d3",x"c0"),
  2288 => (x"e1",x"ca",x"49",x"e0"),
  2289 => (x"de",x"d9",x"c2",x"87"),
  2290 => (x"87",x"c6",x"c0",x"58"),
  2291 => (x"48",x"da",x"d9",x"c2"),
  2292 => (x"49",x"74",x"78",x"c0"),
  2293 => (x"c0",x"05",x"99",x"c2"),
  2294 => (x"eb",x"c3",x"87",x"ce"),
  2295 => (x"87",x"f8",x"e0",x"49"),
  2296 => (x"99",x"c2",x"49",x"70"),
  2297 => (x"87",x"ce",x"c0",x"02"),
  2298 => (x"4a",x"a5",x"d8",x"c1"),
  2299 => (x"c5",x"c0",x"02",x"6a"),
  2300 => (x"49",x"fb",x"4b",x"87"),
  2301 => (x"49",x"74",x"0f",x"73"),
  2302 => (x"c0",x"05",x"99",x"c1"),
  2303 => (x"f4",x"c3",x"87",x"ce"),
  2304 => (x"87",x"d4",x"e0",x"49"),
  2305 => (x"99",x"c2",x"49",x"70"),
  2306 => (x"87",x"cf",x"c0",x"02"),
  2307 => (x"7e",x"a5",x"d8",x"c1"),
  2308 => (x"c0",x"02",x"bf",x"6e"),
  2309 => (x"fa",x"4b",x"87",x"c5"),
  2310 => (x"74",x"0f",x"73",x"49"),
  2311 => (x"05",x"99",x"c8",x"49"),
  2312 => (x"c3",x"87",x"cf",x"c0"),
  2313 => (x"df",x"ff",x"49",x"f5"),
  2314 => (x"49",x"70",x"87",x"ee"),
  2315 => (x"c0",x"02",x"99",x"c2"),
  2316 => (x"f9",x"c2",x"87",x"e6"),
  2317 => (x"c0",x"02",x"bf",x"e1"),
  2318 => (x"c1",x"48",x"87",x"ca"),
  2319 => (x"e5",x"f9",x"c2",x"88"),
  2320 => (x"87",x"cf",x"c0",x"58"),
  2321 => (x"7e",x"a5",x"d8",x"c1"),
  2322 => (x"c0",x"02",x"bf",x"6e"),
  2323 => (x"ff",x"4b",x"87",x"c5"),
  2324 => (x"c4",x"0f",x"73",x"49"),
  2325 => (x"78",x"c1",x"48",x"a6"),
  2326 => (x"99",x"c4",x"49",x"74"),
  2327 => (x"87",x"cf",x"c0",x"05"),
  2328 => (x"ff",x"49",x"f2",x"c3"),
  2329 => (x"70",x"87",x"f1",x"de"),
  2330 => (x"02",x"99",x"c2",x"49"),
  2331 => (x"c2",x"87",x"ec",x"c0"),
  2332 => (x"7e",x"bf",x"e1",x"f9"),
  2333 => (x"a8",x"b7",x"c7",x"48"),
  2334 => (x"87",x"cb",x"c0",x"03"),
  2335 => (x"80",x"c1",x"48",x"6e"),
  2336 => (x"58",x"e5",x"f9",x"c2"),
  2337 => (x"c1",x"87",x"cf",x"c0"),
  2338 => (x"6e",x"7e",x"a5",x"d8"),
  2339 => (x"c5",x"c0",x"02",x"bf"),
  2340 => (x"49",x"fe",x"4b",x"87"),
  2341 => (x"a6",x"c4",x"0f",x"73"),
  2342 => (x"c3",x"78",x"c1",x"48"),
  2343 => (x"dd",x"ff",x"49",x"fd"),
  2344 => (x"49",x"70",x"87",x"f6"),
  2345 => (x"c0",x"02",x"99",x"c2"),
  2346 => (x"f9",x"c2",x"87",x"e5"),
  2347 => (x"c0",x"02",x"bf",x"e1"),
  2348 => (x"f9",x"c2",x"87",x"c9"),
  2349 => (x"78",x"c0",x"48",x"e1"),
  2350 => (x"c1",x"87",x"cf",x"c0"),
  2351 => (x"6e",x"7e",x"a5",x"d8"),
  2352 => (x"c5",x"c0",x"02",x"bf"),
  2353 => (x"49",x"fd",x"4b",x"87"),
  2354 => (x"a6",x"c4",x"0f",x"73"),
  2355 => (x"c3",x"78",x"c1",x"48"),
  2356 => (x"dd",x"ff",x"49",x"fa"),
  2357 => (x"49",x"70",x"87",x"c2"),
  2358 => (x"c0",x"02",x"99",x"c2"),
  2359 => (x"f9",x"c2",x"87",x"e9"),
  2360 => (x"c7",x"48",x"bf",x"e1"),
  2361 => (x"c0",x"03",x"a8",x"b7"),
  2362 => (x"f9",x"c2",x"87",x"c9"),
  2363 => (x"78",x"c7",x"48",x"e1"),
  2364 => (x"c1",x"87",x"cf",x"c0"),
  2365 => (x"6e",x"7e",x"a5",x"d8"),
  2366 => (x"c5",x"c0",x"02",x"bf"),
  2367 => (x"49",x"fc",x"4b",x"87"),
  2368 => (x"a6",x"c4",x"0f",x"73"),
  2369 => (x"c0",x"78",x"c1",x"48"),
  2370 => (x"dc",x"f9",x"c2",x"4b"),
  2371 => (x"cb",x"50",x"c0",x"48"),
  2372 => (x"d1",x"c5",x"49",x"ee"),
  2373 => (x"58",x"a6",x"cc",x"87"),
  2374 => (x"97",x"dc",x"f9",x"c2"),
  2375 => (x"de",x"c1",x"05",x"bf"),
  2376 => (x"c3",x"49",x"74",x"87"),
  2377 => (x"c0",x"05",x"99",x"f0"),
  2378 => (x"da",x"c1",x"87",x"cd"),
  2379 => (x"e7",x"db",x"ff",x"49"),
  2380 => (x"02",x"98",x"70",x"87"),
  2381 => (x"c1",x"87",x"c8",x"c1"),
  2382 => (x"4c",x"bf",x"e8",x"4b"),
  2383 => (x"99",x"ff",x"c3",x"49"),
  2384 => (x"71",x"2c",x"b7",x"c8"),
  2385 => (x"de",x"d9",x"c2",x"b4"),
  2386 => (x"d8",x"ff",x"49",x"bf"),
  2387 => (x"66",x"c8",x"87",x"c0"),
  2388 => (x"87",x"de",x"c4",x"49"),
  2389 => (x"c0",x"02",x"98",x"70"),
  2390 => (x"f9",x"c2",x"87",x"c6"),
  2391 => (x"50",x"c1",x"48",x"dc"),
  2392 => (x"97",x"dc",x"f9",x"c2"),
  2393 => (x"d6",x"c0",x"05",x"bf"),
  2394 => (x"c3",x"49",x"74",x"87"),
  2395 => (x"ff",x"05",x"99",x"f0"),
  2396 => (x"da",x"c1",x"87",x"c5"),
  2397 => (x"df",x"da",x"ff",x"49"),
  2398 => (x"05",x"98",x"70",x"87"),
  2399 => (x"73",x"87",x"f8",x"fe"),
  2400 => (x"dc",x"c0",x"02",x"9b"),
  2401 => (x"48",x"a6",x"c8",x"87"),
  2402 => (x"bf",x"e1",x"f9",x"c2"),
  2403 => (x"49",x"66",x"c8",x"78"),
  2404 => (x"a1",x"75",x"91",x"cb"),
  2405 => (x"02",x"bf",x"6e",x"7e"),
  2406 => (x"4b",x"87",x"c6",x"c0"),
  2407 => (x"73",x"49",x"66",x"c8"),
  2408 => (x"02",x"66",x"c4",x"0f"),
  2409 => (x"c2",x"87",x"c8",x"c0"),
  2410 => (x"49",x"bf",x"e1",x"f9"),
  2411 => (x"c2",x"87",x"f8",x"ee"),
  2412 => (x"02",x"bf",x"e2",x"d9"),
  2413 => (x"49",x"87",x"dd",x"c0"),
  2414 => (x"70",x"87",x"f7",x"c2"),
  2415 => (x"d3",x"c0",x"02",x"98"),
  2416 => (x"e1",x"f9",x"c2",x"87"),
  2417 => (x"de",x"ee",x"49",x"bf"),
  2418 => (x"ef",x"49",x"c0",x"87"),
  2419 => (x"d9",x"c2",x"87",x"fe"),
  2420 => (x"78",x"c0",x"48",x"e2"),
  2421 => (x"d8",x"ef",x"8e",x"f4"),
  2422 => (x"79",x"6f",x"4a",x"87"),
  2423 => (x"73",x"79",x"65",x"6b"),
  2424 => (x"00",x"6e",x"6f",x"20"),
  2425 => (x"6b",x"79",x"6f",x"4a"),
  2426 => (x"20",x"73",x"79",x"65"),
  2427 => (x"00",x"66",x"66",x"6f"),
  2428 => (x"5c",x"5b",x"5e",x"0e"),
  2429 => (x"71",x"1e",x"0e",x"5d"),
  2430 => (x"dd",x"f9",x"c2",x"4c"),
  2431 => (x"cd",x"c1",x"49",x"bf"),
  2432 => (x"d1",x"c1",x"4d",x"a1"),
  2433 => (x"74",x"7e",x"69",x"81"),
  2434 => (x"87",x"cf",x"02",x"9c"),
  2435 => (x"74",x"4b",x"a5",x"c4"),
  2436 => (x"dd",x"f9",x"c2",x"7b"),
  2437 => (x"e0",x"ee",x"49",x"bf"),
  2438 => (x"74",x"7b",x"6e",x"87"),
  2439 => (x"87",x"c4",x"05",x"9c"),
  2440 => (x"87",x"c2",x"4b",x"c0"),
  2441 => (x"49",x"73",x"4b",x"c1"),
  2442 => (x"d4",x"87",x"e1",x"ee"),
  2443 => (x"87",x"c8",x"02",x"66"),
  2444 => (x"87",x"f2",x"c0",x"49"),
  2445 => (x"87",x"c2",x"4a",x"70"),
  2446 => (x"d9",x"c2",x"4a",x"c0"),
  2447 => (x"ed",x"26",x"5a",x"e6"),
  2448 => (x"00",x"00",x"87",x"ef"),
  2449 => (x"00",x"00",x"00",x"00"),
  2450 => (x"12",x"58",x"00",x"00"),
  2451 => (x"1b",x"1d",x"14",x"11"),
  2452 => (x"59",x"5a",x"23",x"1c"),
  2453 => (x"f2",x"f5",x"94",x"91"),
  2454 => (x"00",x"00",x"f4",x"eb"),
  2455 => (x"00",x"00",x"00",x"00"),
  2456 => (x"00",x"00",x"00",x"00"),
  2457 => (x"71",x"1e",x"00",x"00"),
  2458 => (x"bf",x"c8",x"ff",x"4a"),
  2459 => (x"48",x"a1",x"72",x"49"),
  2460 => (x"ff",x"1e",x"4f",x"26"),
  2461 => (x"fe",x"89",x"bf",x"c8"),
  2462 => (x"c0",x"c0",x"c0",x"c0"),
  2463 => (x"c4",x"01",x"a9",x"c0"),
  2464 => (x"c2",x"4a",x"c0",x"87"),
  2465 => (x"72",x"4a",x"c1",x"87"),
  2466 => (x"0e",x"4f",x"26",x"48"),
  2467 => (x"5d",x"5c",x"5b",x"5e"),
  2468 => (x"ff",x"4b",x"71",x"0e"),
  2469 => (x"66",x"d0",x"4c",x"d4"),
  2470 => (x"d6",x"78",x"c0",x"48"),
  2471 => (x"ef",x"d7",x"ff",x"49"),
  2472 => (x"7c",x"ff",x"c3",x"87"),
  2473 => (x"ff",x"c3",x"49",x"6c"),
  2474 => (x"49",x"4d",x"71",x"99"),
  2475 => (x"c1",x"99",x"f0",x"c3"),
  2476 => (x"cb",x"05",x"a9",x"e0"),
  2477 => (x"7c",x"ff",x"c3",x"87"),
  2478 => (x"98",x"c3",x"48",x"6c"),
  2479 => (x"78",x"08",x"66",x"d0"),
  2480 => (x"6c",x"7c",x"ff",x"c3"),
  2481 => (x"31",x"c8",x"49",x"4a"),
  2482 => (x"6c",x"7c",x"ff",x"c3"),
  2483 => (x"72",x"b2",x"71",x"4a"),
  2484 => (x"c3",x"31",x"c8",x"49"),
  2485 => (x"4a",x"6c",x"7c",x"ff"),
  2486 => (x"49",x"72",x"b2",x"71"),
  2487 => (x"ff",x"c3",x"31",x"c8"),
  2488 => (x"71",x"4a",x"6c",x"7c"),
  2489 => (x"48",x"d0",x"ff",x"b2"),
  2490 => (x"73",x"78",x"e0",x"c0"),
  2491 => (x"87",x"c2",x"02",x"9b"),
  2492 => (x"48",x"75",x"7b",x"72"),
  2493 => (x"4c",x"26",x"4d",x"26"),
  2494 => (x"4f",x"26",x"4b",x"26"),
  2495 => (x"0e",x"4f",x"26",x"1e"),
  2496 => (x"0e",x"5c",x"5b",x"5e"),
  2497 => (x"1e",x"76",x"86",x"f8"),
  2498 => (x"fd",x"49",x"a6",x"c8"),
  2499 => (x"86",x"c4",x"87",x"fd"),
  2500 => (x"48",x"6e",x"4b",x"70"),
  2501 => (x"c2",x"03",x"a8",x"c2"),
  2502 => (x"4a",x"73",x"87",x"f0"),
  2503 => (x"c1",x"9a",x"f0",x"c3"),
  2504 => (x"c7",x"02",x"aa",x"d0"),
  2505 => (x"aa",x"e0",x"c1",x"87"),
  2506 => (x"87",x"de",x"c2",x"05"),
  2507 => (x"99",x"c8",x"49",x"73"),
  2508 => (x"ff",x"87",x"c3",x"02"),
  2509 => (x"4c",x"73",x"87",x"c6"),
  2510 => (x"ac",x"c2",x"9c",x"c3"),
  2511 => (x"87",x"c2",x"c1",x"05"),
  2512 => (x"c9",x"49",x"66",x"c4"),
  2513 => (x"c4",x"1e",x"71",x"31"),
  2514 => (x"92",x"d4",x"4a",x"66"),
  2515 => (x"49",x"e5",x"f9",x"c2"),
  2516 => (x"c9",x"fe",x"81",x"72"),
  2517 => (x"49",x"d8",x"87",x"f1"),
  2518 => (x"87",x"f4",x"d4",x"ff"),
  2519 => (x"c2",x"1e",x"c0",x"c8"),
  2520 => (x"fd",x"49",x"ce",x"e8"),
  2521 => (x"ff",x"87",x"f7",x"e5"),
  2522 => (x"e0",x"c0",x"48",x"d0"),
  2523 => (x"ce",x"e8",x"c2",x"78"),
  2524 => (x"4a",x"66",x"cc",x"1e"),
  2525 => (x"f9",x"c2",x"92",x"d4"),
  2526 => (x"81",x"72",x"49",x"e5"),
  2527 => (x"87",x"f9",x"c7",x"fe"),
  2528 => (x"ac",x"c1",x"86",x"cc"),
  2529 => (x"87",x"c2",x"c1",x"05"),
  2530 => (x"c9",x"49",x"66",x"c4"),
  2531 => (x"c4",x"1e",x"71",x"31"),
  2532 => (x"92",x"d4",x"4a",x"66"),
  2533 => (x"49",x"e5",x"f9",x"c2"),
  2534 => (x"c8",x"fe",x"81",x"72"),
  2535 => (x"e8",x"c2",x"87",x"e9"),
  2536 => (x"66",x"c8",x"1e",x"ce"),
  2537 => (x"c2",x"92",x"d4",x"4a"),
  2538 => (x"72",x"49",x"e5",x"f9"),
  2539 => (x"fa",x"c5",x"fe",x"81"),
  2540 => (x"ff",x"49",x"d7",x"87"),
  2541 => (x"c8",x"87",x"d9",x"d3"),
  2542 => (x"e8",x"c2",x"1e",x"c0"),
  2543 => (x"e3",x"fd",x"49",x"ce"),
  2544 => (x"86",x"cc",x"87",x"f5"),
  2545 => (x"c0",x"48",x"d0",x"ff"),
  2546 => (x"8e",x"f8",x"78",x"e0"),
  2547 => (x"0e",x"87",x"e7",x"fc"),
  2548 => (x"5d",x"5c",x"5b",x"5e"),
  2549 => (x"ff",x"4a",x"71",x"0e"),
  2550 => (x"66",x"d0",x"4c",x"d4"),
  2551 => (x"ad",x"b7",x"c3",x"4d"),
  2552 => (x"c0",x"87",x"c5",x"06"),
  2553 => (x"87",x"e1",x"c1",x"48"),
  2554 => (x"4b",x"75",x"1e",x"72"),
  2555 => (x"f9",x"c2",x"93",x"d4"),
  2556 => (x"49",x"73",x"83",x"e5"),
  2557 => (x"87",x"c1",x"c0",x"fe"),
  2558 => (x"4b",x"6b",x"83",x"c8"),
  2559 => (x"c8",x"48",x"d0",x"ff"),
  2560 => (x"7c",x"dd",x"78",x"e1"),
  2561 => (x"ff",x"c3",x"48",x"73"),
  2562 => (x"73",x"7c",x"70",x"98"),
  2563 => (x"29",x"b7",x"c8",x"49"),
  2564 => (x"ff",x"c3",x"48",x"71"),
  2565 => (x"73",x"7c",x"70",x"98"),
  2566 => (x"29",x"b7",x"d0",x"49"),
  2567 => (x"ff",x"c3",x"48",x"71"),
  2568 => (x"73",x"7c",x"70",x"98"),
  2569 => (x"28",x"b7",x"d8",x"48"),
  2570 => (x"7c",x"c0",x"7c",x"70"),
  2571 => (x"7c",x"7c",x"7c",x"7c"),
  2572 => (x"7c",x"7c",x"7c",x"7c"),
  2573 => (x"ff",x"7c",x"7c",x"7c"),
  2574 => (x"e0",x"c0",x"48",x"d0"),
  2575 => (x"dc",x"1e",x"75",x"78"),
  2576 => (x"f0",x"d1",x"ff",x"49"),
  2577 => (x"73",x"86",x"c8",x"87"),
  2578 => (x"87",x"e8",x"fa",x"48"),
  2579 => (x"c4",x"4a",x"71",x"1e"),
  2580 => (x"f9",x"c2",x"49",x"a2"),
  2581 => (x"78",x"6a",x"48",x"c8"),
  2582 => (x"48",x"c2",x"d9",x"c2"),
  2583 => (x"d9",x"c2",x"78",x"69"),
  2584 => (x"e6",x"49",x"bf",x"c2"),
  2585 => (x"d1",x"ff",x"87",x"f4"),
  2586 => (x"4f",x"26",x"87",x"fd"),
  2587 => (x"c4",x"4a",x"71",x"1e"),
  2588 => (x"f9",x"c2",x"49",x"a2"),
  2589 => (x"c2",x"7a",x"bf",x"c8"),
  2590 => (x"79",x"bf",x"c2",x"d9"),
  2591 => (x"71",x"1e",x"4f",x"26"),
  2592 => (x"c0",x"02",x"9a",x"4a"),
  2593 => (x"c2",x"1e",x"87",x"ee"),
  2594 => (x"fd",x"49",x"c4",x"f5"),
  2595 => (x"c4",x"87",x"ea",x"fd"),
  2596 => (x"02",x"98",x"70",x"86"),
  2597 => (x"e8",x"c2",x"87",x"de"),
  2598 => (x"f5",x"c2",x"1e",x"ce"),
  2599 => (x"c2",x"fe",x"49",x"c4"),
  2600 => (x"86",x"c4",x"87",x"c9"),
  2601 => (x"cb",x"02",x"98",x"70"),
  2602 => (x"ce",x"e8",x"c2",x"87"),
  2603 => (x"87",x"dc",x"fe",x"49"),
  2604 => (x"87",x"c2",x"48",x"c1"),
  2605 => (x"4f",x"26",x"48",x"c0"),
  2606 => (x"9a",x"4a",x"71",x"1e"),
  2607 => (x"87",x"ee",x"c0",x"02"),
  2608 => (x"c4",x"f5",x"c2",x"1e"),
  2609 => (x"f0",x"fc",x"fd",x"49"),
  2610 => (x"70",x"86",x"c4",x"87"),
  2611 => (x"87",x"de",x"02",x"98"),
  2612 => (x"49",x"ce",x"e8",x"c2"),
  2613 => (x"c2",x"87",x"d5",x"fe"),
  2614 => (x"c2",x"1e",x"ce",x"e8"),
  2615 => (x"fe",x"49",x"c4",x"f5"),
  2616 => (x"c4",x"87",x"d6",x"c2"),
  2617 => (x"02",x"98",x"70",x"86"),
  2618 => (x"48",x"c1",x"87",x"c4"),
  2619 => (x"48",x"c0",x"87",x"c2"),
  2620 => (x"c1",x"1e",x"4f",x"26"),
  2621 => (x"c0",x"48",x"cc",x"e7"),
  2622 => (x"cd",x"fa",x"c2",x"50"),
  2623 => (x"87",x"cc",x"05",x"bf"),
  2624 => (x"49",x"ff",x"e4",x"c2"),
  2625 => (x"87",x"e1",x"d5",x"fe"),
  2626 => (x"58",x"d1",x"fa",x"c2"),
  2627 => (x"48",x"cc",x"e7",x"c1"),
  2628 => (x"fa",x"c2",x"50",x"c2"),
  2629 => (x"cc",x"05",x"bf",x"d1"),
  2630 => (x"cb",x"e5",x"c2",x"87"),
  2631 => (x"c8",x"d5",x"fe",x"49"),
  2632 => (x"d5",x"fa",x"c2",x"87"),
  2633 => (x"d5",x"fa",x"c2",x"58"),
  2634 => (x"87",x"d1",x"05",x"bf"),
  2635 => (x"c2",x"1e",x"f1",x"c0"),
  2636 => (x"fe",x"49",x"d7",x"e5"),
  2637 => (x"c4",x"87",x"c5",x"db"),
  2638 => (x"d9",x"fa",x"c2",x"86"),
  2639 => (x"56",x"4f",x"26",x"58"),
  2640 => (x"30",x"32",x"43",x"49"),
  2641 => (x"52",x"20",x"20",x"20"),
  2642 => (x"4d",x"00",x"4d",x"4f"),
  2643 => (x"43",x"41",x"47",x"45"),
  2644 => (x"52",x"54",x"52",x"41"),
  2645 => (x"4d",x"00",x"4d",x"4f"),
  2646 => (x"43",x"41",x"47",x"45"),
  2647 => (x"4e",x"54",x"52",x"41"),
  2648 => (x"1e",x"00",x"20",x"56"),
  2649 => (x"4b",x"c0",x"1e",x"73"),
  2650 => (x"48",x"cd",x"fa",x"c2"),
  2651 => (x"fa",x"c2",x"78",x"c0"),
  2652 => (x"78",x"c0",x"48",x"d1"),
  2653 => (x"48",x"d5",x"fa",x"c2"),
  2654 => (x"f5",x"fd",x"78",x"c0"),
  2655 => (x"d1",x"e7",x"c2",x"87"),
  2656 => (x"c4",x"f5",x"c2",x"1e"),
  2657 => (x"f0",x"f9",x"fd",x"49"),
  2658 => (x"70",x"86",x"c4",x"87"),
  2659 => (x"87",x"c9",x"02",x"98"),
  2660 => (x"bf",x"c8",x"f5",x"c2"),
  2661 => (x"d0",x"c2",x"fe",x"49"),
  2662 => (x"87",x"d6",x"fd",x"87"),
  2663 => (x"c2",x"fe",x"49",x"c0"),
  2664 => (x"fa",x"c2",x"87",x"c7"),
  2665 => (x"cd",x"02",x"bf",x"d1"),
  2666 => (x"c8",x"f9",x"c2",x"87"),
  2667 => (x"c0",x"c8",x"48",x"bf"),
  2668 => (x"f9",x"c2",x"b0",x"c0"),
  2669 => (x"cc",x"ff",x"58",x"cc"),
  2670 => (x"fa",x"c2",x"87",x"ed"),
  2671 => (x"c4",x"05",x"bf",x"cd"),
  2672 => (x"dd",x"e7",x"c2",x"87"),
  2673 => (x"c4",x"48",x"73",x"4b"),
  2674 => (x"26",x"4d",x"26",x"87"),
  2675 => (x"26",x"4b",x"26",x"4c"),
  2676 => (x"41",x"48",x"43",x"4f"),
  2677 => (x"20",x"30",x"32",x"4d"),
  2678 => (x"20",x"20",x"20",x"20"),
  2679 => (x"4d",x"4f",x"52",x"00"),
  2680 => (x"69",x"61",x"66",x"20"),
  2681 => (x"00",x"64",x"65",x"6c"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

